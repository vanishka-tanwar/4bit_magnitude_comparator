magic
tech sky130A
magscale 1 2
timestamp 1629539722
<< checkpaint >>
rect -3932 -3932 12662 14806
<< viali >>
rect 4445 8041 4479 8075
rect 1777 7973 1811 8007
rect 1961 7837 1995 7871
rect 6837 7837 6871 7871
rect 4537 7769 4571 7803
rect 6653 7701 6687 7735
rect 1409 7361 1443 7395
rect 6837 7361 6871 7395
rect 1593 7157 1627 7191
rect 6653 7157 6687 7191
rect 4445 5865 4479 5899
rect 3985 5661 4019 5695
rect 4445 5661 4479 5695
rect 4629 5661 4663 5695
rect 5457 5661 5491 5695
rect 3893 5525 3927 5559
rect 5365 5525 5399 5559
rect 5365 5321 5399 5355
rect 6469 5253 6503 5287
rect 3433 5185 3467 5219
rect 3617 5185 3651 5219
rect 4077 5185 4111 5219
rect 4721 5185 4755 5219
rect 4900 5185 4934 5219
rect 5000 5185 5034 5219
rect 5089 5185 5123 5219
rect 6377 5185 6411 5219
rect 3617 4981 3651 5015
rect 4169 4981 4203 5015
rect 4261 4777 4295 4811
rect 4905 4777 4939 4811
rect 1593 4709 1627 4743
rect 3065 4641 3099 4675
rect 5365 4641 5399 4675
rect 1409 4573 1443 4607
rect 3193 4573 3227 4607
rect 3985 4573 4019 4607
rect 4077 4573 4111 4607
rect 4353 4573 4387 4607
rect 5089 4573 5123 4607
rect 5273 4573 5307 4607
rect 5457 4573 5491 4607
rect 5641 4573 5675 4607
rect 2789 4505 2823 4539
rect 2973 4505 3007 4539
rect 3065 4505 3099 4539
rect 6653 4505 6687 4539
rect 3801 4437 3835 4471
rect 6745 4437 6779 4471
rect 3801 4233 3835 4267
rect 4721 4233 4755 4267
rect 3065 4097 3099 4131
rect 3249 4097 3283 4131
rect 3617 4097 3651 4131
rect 4905 4097 4939 4131
rect 5181 4097 5215 4131
rect 5365 4097 5399 4131
rect 3341 4029 3375 4063
rect 3433 4029 3467 4063
rect 3893 3689 3927 3723
rect 5089 3689 5123 3723
rect 3801 3485 3835 3519
rect 4997 3485 5031 3519
rect 5191 3485 5225 3519
rect 5825 3485 5859 3519
rect 5733 3417 5767 3451
rect 1593 2601 1627 2635
rect 3249 2601 3283 2635
rect 5641 2601 5675 2635
rect 6653 2601 6687 2635
rect 1409 2397 1443 2431
rect 3065 2397 3099 2431
rect 5825 2397 5859 2431
rect 6837 2397 6871 2431
<< metal1 >>
rect 1104 8186 7544 8208
rect 1104 8134 2055 8186
rect 2107 8134 2119 8186
rect 2171 8134 2183 8186
rect 2235 8134 2247 8186
rect 2299 8134 4202 8186
rect 4254 8134 4266 8186
rect 4318 8134 4330 8186
rect 4382 8134 4394 8186
rect 4446 8134 6348 8186
rect 6400 8134 6412 8186
rect 6464 8134 6476 8186
rect 6528 8134 6540 8186
rect 6592 8134 7544 8186
rect 1104 8112 7544 8134
rect 4433 8075 4491 8081
rect 4433 8041 4445 8075
rect 4479 8072 4491 8075
rect 4522 8072 4528 8084
rect 4479 8044 4528 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 4522 8032 4528 8044
rect 4580 8032 4586 8084
rect 1302 7964 1308 8016
rect 1360 8004 1366 8016
rect 1765 8007 1823 8013
rect 1765 8004 1777 8007
rect 1360 7976 1777 8004
rect 1360 7964 1366 7976
rect 1765 7973 1777 7976
rect 1811 7973 1823 8007
rect 1765 7967 1823 7973
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7868 2007 7871
rect 4614 7868 4620 7880
rect 1995 7840 4620 7868
rect 1995 7837 2007 7840
rect 1949 7831 2007 7837
rect 4614 7828 4620 7840
rect 4672 7828 4678 7880
rect 6825 7871 6883 7877
rect 6825 7837 6837 7871
rect 6871 7868 6883 7871
rect 7190 7868 7196 7880
rect 6871 7840 7196 7868
rect 6871 7837 6883 7840
rect 6825 7831 6883 7837
rect 7190 7828 7196 7840
rect 7248 7828 7254 7880
rect 4522 7800 4528 7812
rect 4483 7772 4528 7800
rect 4522 7760 4528 7772
rect 4580 7760 4586 7812
rect 5626 7692 5632 7744
rect 5684 7732 5690 7744
rect 6641 7735 6699 7741
rect 6641 7732 6653 7735
rect 5684 7704 6653 7732
rect 5684 7692 5690 7704
rect 6641 7701 6653 7704
rect 6687 7701 6699 7735
rect 6641 7695 6699 7701
rect 1104 7642 7544 7664
rect 1104 7590 3128 7642
rect 3180 7590 3192 7642
rect 3244 7590 3256 7642
rect 3308 7590 3320 7642
rect 3372 7590 5275 7642
rect 5327 7590 5339 7642
rect 5391 7590 5403 7642
rect 5455 7590 5467 7642
rect 5519 7590 7544 7642
rect 1104 7568 7544 7590
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 6822 7392 6828 7404
rect 6783 7364 6828 7392
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 1581 7191 1639 7197
rect 1581 7157 1593 7191
rect 1627 7188 1639 7191
rect 4798 7188 4804 7200
rect 1627 7160 4804 7188
rect 1627 7157 1639 7160
rect 1581 7151 1639 7157
rect 4798 7148 4804 7160
rect 4856 7148 4862 7200
rect 6638 7188 6644 7200
rect 6599 7160 6644 7188
rect 6638 7148 6644 7160
rect 6696 7148 6702 7200
rect 1104 7098 7544 7120
rect 1104 7046 2055 7098
rect 2107 7046 2119 7098
rect 2171 7046 2183 7098
rect 2235 7046 2247 7098
rect 2299 7046 4202 7098
rect 4254 7046 4266 7098
rect 4318 7046 4330 7098
rect 4382 7046 4394 7098
rect 4446 7046 6348 7098
rect 6400 7046 6412 7098
rect 6464 7046 6476 7098
rect 6528 7046 6540 7098
rect 6592 7046 7544 7098
rect 1104 7024 7544 7046
rect 1104 6554 7544 6576
rect 1104 6502 3128 6554
rect 3180 6502 3192 6554
rect 3244 6502 3256 6554
rect 3308 6502 3320 6554
rect 3372 6502 5275 6554
rect 5327 6502 5339 6554
rect 5391 6502 5403 6554
rect 5455 6502 5467 6554
rect 5519 6502 7544 6554
rect 1104 6480 7544 6502
rect 1104 6010 7544 6032
rect 1104 5958 2055 6010
rect 2107 5958 2119 6010
rect 2171 5958 2183 6010
rect 2235 5958 2247 6010
rect 2299 5958 4202 6010
rect 4254 5958 4266 6010
rect 4318 5958 4330 6010
rect 4382 5958 4394 6010
rect 4446 5958 6348 6010
rect 6400 5958 6412 6010
rect 6464 5958 6476 6010
rect 6528 5958 6540 6010
rect 6592 5958 7544 6010
rect 1104 5936 7544 5958
rect 4433 5899 4491 5905
rect 4433 5865 4445 5899
rect 4479 5896 4491 5899
rect 4522 5896 4528 5908
rect 4479 5868 4528 5896
rect 4479 5865 4491 5868
rect 4433 5859 4491 5865
rect 4522 5856 4528 5868
rect 4580 5856 4586 5908
rect 6638 5760 6644 5772
rect 3988 5732 6644 5760
rect 3988 5701 4016 5732
rect 6638 5720 6644 5732
rect 6696 5720 6702 5772
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4522 5692 4528 5704
rect 4479 5664 4528 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 4614 5652 4620 5704
rect 4672 5692 4678 5704
rect 4672 5664 4717 5692
rect 4672 5652 4678 5664
rect 4982 5652 4988 5704
rect 5040 5692 5046 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5040 5664 5457 5692
rect 5040 5652 5046 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 3418 5516 3424 5568
rect 3476 5556 3482 5568
rect 3881 5559 3939 5565
rect 3881 5556 3893 5559
rect 3476 5528 3893 5556
rect 3476 5516 3482 5528
rect 3881 5525 3893 5528
rect 3927 5525 3939 5559
rect 3881 5519 3939 5525
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 5353 5559 5411 5565
rect 5353 5556 5365 5559
rect 5224 5528 5365 5556
rect 5224 5516 5230 5528
rect 5353 5525 5365 5528
rect 5399 5525 5411 5559
rect 5353 5519 5411 5525
rect 1104 5466 7544 5488
rect 1104 5414 3128 5466
rect 3180 5414 3192 5466
rect 3244 5414 3256 5466
rect 3308 5414 3320 5466
rect 3372 5414 5275 5466
rect 5327 5414 5339 5466
rect 5391 5414 5403 5466
rect 5455 5414 5467 5466
rect 5519 5414 7544 5466
rect 1104 5392 7544 5414
rect 4522 5312 4528 5364
rect 4580 5352 4586 5364
rect 5353 5355 5411 5361
rect 5353 5352 5365 5355
rect 4580 5324 5365 5352
rect 4580 5312 4586 5324
rect 5353 5321 5365 5324
rect 5399 5321 5411 5355
rect 5353 5315 5411 5321
rect 6457 5287 6515 5293
rect 6457 5284 6469 5287
rect 5092 5256 6469 5284
rect 3421 5219 3479 5225
rect 3421 5185 3433 5219
rect 3467 5185 3479 5219
rect 3602 5216 3608 5228
rect 3563 5188 3608 5216
rect 3421 5179 3479 5185
rect 3050 5108 3056 5160
rect 3108 5148 3114 5160
rect 3436 5148 3464 5179
rect 3602 5176 3608 5188
rect 3660 5176 3666 5228
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 4890 5225 4896 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 3844 5188 4077 5216
rect 3844 5176 3850 5188
rect 4065 5185 4077 5188
rect 4111 5216 4123 5219
rect 4709 5219 4767 5225
rect 4709 5216 4721 5219
rect 4111 5188 4721 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4709 5185 4721 5188
rect 4755 5185 4767 5219
rect 4888 5216 4896 5225
rect 4851 5188 4896 5216
rect 4709 5179 4767 5185
rect 4888 5179 4896 5188
rect 4890 5176 4896 5179
rect 4948 5176 4954 5228
rect 5092 5225 5120 5256
rect 6457 5253 6469 5256
rect 6503 5253 6515 5287
rect 6457 5247 6515 5253
rect 4988 5219 5046 5225
rect 4988 5185 5000 5219
rect 5034 5185 5046 5219
rect 4988 5179 5046 5185
rect 5077 5219 5135 5225
rect 5077 5185 5089 5219
rect 5123 5185 5135 5219
rect 5077 5179 5135 5185
rect 3108 5120 4660 5148
rect 3108 5108 3114 5120
rect 3605 5015 3663 5021
rect 3605 4981 3617 5015
rect 3651 5012 3663 5015
rect 4062 5012 4068 5024
rect 3651 4984 4068 5012
rect 3651 4981 3663 4984
rect 3605 4975 3663 4981
rect 4062 4972 4068 4984
rect 4120 4972 4126 5024
rect 4157 5015 4215 5021
rect 4157 4981 4169 5015
rect 4203 5012 4215 5015
rect 4522 5012 4528 5024
rect 4203 4984 4528 5012
rect 4203 4981 4215 4984
rect 4157 4975 4215 4981
rect 4522 4972 4528 4984
rect 4580 4972 4586 5024
rect 4632 5012 4660 5120
rect 5003 5092 5031 5179
rect 5442 5176 5448 5228
rect 5500 5216 5506 5228
rect 6365 5219 6423 5225
rect 6365 5216 6377 5219
rect 5500 5188 6377 5216
rect 5500 5176 5506 5188
rect 6365 5185 6377 5188
rect 6411 5185 6423 5219
rect 6365 5179 6423 5185
rect 4982 5040 4988 5092
rect 5040 5040 5046 5092
rect 5626 5012 5632 5024
rect 4632 4984 5632 5012
rect 5626 4972 5632 4984
rect 5684 4972 5690 5024
rect 1104 4922 7544 4944
rect 1104 4870 2055 4922
rect 2107 4870 2119 4922
rect 2171 4870 2183 4922
rect 2235 4870 2247 4922
rect 2299 4870 4202 4922
rect 4254 4870 4266 4922
rect 4318 4870 4330 4922
rect 4382 4870 4394 4922
rect 4446 4870 6348 4922
rect 6400 4870 6412 4922
rect 6464 4870 6476 4922
rect 6528 4870 6540 4922
rect 6592 4870 7544 4922
rect 1104 4848 7544 4870
rect 4249 4811 4307 4817
rect 4249 4777 4261 4811
rect 4295 4808 4307 4811
rect 4522 4808 4528 4820
rect 4295 4780 4528 4808
rect 4295 4777 4307 4780
rect 4249 4771 4307 4777
rect 4522 4768 4528 4780
rect 4580 4768 4586 4820
rect 4890 4808 4896 4820
rect 4851 4780 4896 4808
rect 4890 4768 4896 4780
rect 4948 4768 4954 4820
rect 1581 4743 1639 4749
rect 1581 4709 1593 4743
rect 1627 4740 1639 4743
rect 1627 4712 4568 4740
rect 1627 4709 1639 4712
rect 1581 4703 1639 4709
rect 2958 4632 2964 4684
rect 3016 4672 3022 4684
rect 3053 4675 3111 4681
rect 3053 4672 3065 4675
rect 3016 4644 3065 4672
rect 3016 4632 3022 4644
rect 3053 4641 3065 4644
rect 3099 4672 3111 4675
rect 3099 4644 4016 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 1394 4604 1400 4616
rect 1355 4576 1400 4604
rect 1394 4564 1400 4576
rect 1452 4564 1458 4616
rect 3181 4607 3239 4613
rect 3181 4573 3193 4607
rect 3227 4604 3239 4607
rect 3602 4604 3608 4616
rect 3227 4576 3608 4604
rect 3227 4573 3239 4576
rect 3181 4567 3239 4573
rect 3602 4564 3608 4576
rect 3660 4604 3666 4616
rect 3878 4604 3884 4616
rect 3660 4576 3884 4604
rect 3660 4564 3666 4576
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 3988 4613 4016 4644
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 3973 4567 4031 4573
rect 4062 4564 4068 4616
rect 4120 4604 4126 4616
rect 4338 4604 4344 4616
rect 4120 4576 4165 4604
rect 4299 4576 4344 4604
rect 4120 4564 4126 4576
rect 4338 4564 4344 4576
rect 4396 4564 4402 4616
rect 4540 4604 4568 4712
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 5442 4740 5448 4752
rect 4856 4712 5448 4740
rect 4856 4700 4862 4712
rect 5442 4700 5448 4712
rect 5500 4700 5506 4752
rect 5166 4632 5172 4684
rect 5224 4672 5230 4684
rect 5353 4675 5411 4681
rect 5353 4672 5365 4675
rect 5224 4644 5365 4672
rect 5224 4632 5230 4644
rect 5353 4641 5365 4644
rect 5399 4641 5411 4675
rect 5353 4635 5411 4641
rect 5074 4604 5080 4616
rect 4540 4576 5080 4604
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5460 4613 5488 4700
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5445 4607 5503 4613
rect 5445 4573 5457 4607
rect 5491 4573 5503 4607
rect 5626 4604 5632 4616
rect 5587 4576 5632 4604
rect 5445 4567 5503 4573
rect 2774 4496 2780 4548
rect 2832 4536 2838 4548
rect 2961 4539 3019 4545
rect 2832 4508 2877 4536
rect 2832 4496 2838 4508
rect 2961 4505 2973 4539
rect 3007 4505 3019 4539
rect 2961 4499 3019 4505
rect 2976 4468 3004 4499
rect 3050 4496 3056 4548
rect 3108 4536 3114 4548
rect 3510 4536 3516 4548
rect 3108 4508 3516 4536
rect 3108 4496 3114 4508
rect 3510 4496 3516 4508
rect 3568 4496 3574 4548
rect 5166 4496 5172 4548
rect 5224 4536 5230 4548
rect 5276 4536 5304 4567
rect 5626 4564 5632 4576
rect 5684 4564 5690 4616
rect 6641 4539 6699 4545
rect 6641 4536 6653 4539
rect 5224 4508 5304 4536
rect 5368 4508 6653 4536
rect 5224 4496 5230 4508
rect 3418 4468 3424 4480
rect 2976 4440 3424 4468
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 3789 4471 3847 4477
rect 3789 4437 3801 4471
rect 3835 4468 3847 4471
rect 4614 4468 4620 4480
rect 3835 4440 4620 4468
rect 3835 4437 3847 4440
rect 3789 4431 3847 4437
rect 4614 4428 4620 4440
rect 4672 4468 4678 4480
rect 5368 4468 5396 4508
rect 6641 4505 6653 4508
rect 6687 4505 6699 4539
rect 6641 4499 6699 4505
rect 6730 4468 6736 4480
rect 4672 4440 5396 4468
rect 6691 4440 6736 4468
rect 4672 4428 4678 4440
rect 6730 4428 6736 4440
rect 6788 4428 6794 4480
rect 1104 4378 7544 4400
rect 1104 4326 3128 4378
rect 3180 4326 3192 4378
rect 3244 4326 3256 4378
rect 3308 4326 3320 4378
rect 3372 4326 5275 4378
rect 5327 4326 5339 4378
rect 5391 4326 5403 4378
rect 5455 4326 5467 4378
rect 5519 4326 7544 4378
rect 1104 4304 7544 4326
rect 3786 4264 3792 4276
rect 3747 4236 3792 4264
rect 3786 4224 3792 4236
rect 3844 4224 3850 4276
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4709 4267 4767 4273
rect 4709 4264 4721 4267
rect 4396 4236 4721 4264
rect 4396 4224 4402 4236
rect 4709 4233 4721 4236
rect 4755 4233 4767 4267
rect 4709 4227 4767 4233
rect 3418 4196 3424 4208
rect 3252 4168 3424 4196
rect 2958 4088 2964 4140
rect 3016 4128 3022 4140
rect 3252 4137 3280 4168
rect 3418 4156 3424 4168
rect 3476 4156 3482 4208
rect 5074 4156 5080 4208
rect 5132 4196 5138 4208
rect 5132 4168 5396 4196
rect 5132 4156 5138 4168
rect 3053 4131 3111 4137
rect 3053 4128 3065 4131
rect 3016 4100 3065 4128
rect 3016 4088 3022 4100
rect 3053 4097 3065 4100
rect 3099 4097 3111 4131
rect 3053 4091 3111 4097
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3510 4088 3516 4140
rect 3568 4128 3574 4140
rect 3605 4131 3663 4137
rect 3605 4128 3617 4131
rect 3568 4100 3617 4128
rect 3568 4088 3574 4100
rect 3605 4097 3617 4100
rect 3651 4097 3663 4131
rect 4890 4128 4896 4140
rect 4851 4100 4896 4128
rect 3605 4091 3663 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5166 4128 5172 4140
rect 5127 4100 5172 4128
rect 5166 4088 5172 4100
rect 5224 4088 5230 4140
rect 5368 4137 5396 4168
rect 5353 4131 5411 4137
rect 5353 4097 5365 4131
rect 5399 4097 5411 4131
rect 5353 4091 5411 4097
rect 2774 4020 2780 4072
rect 2832 4060 2838 4072
rect 3329 4063 3387 4069
rect 3329 4060 3341 4063
rect 2832 4032 3341 4060
rect 2832 4020 2838 4032
rect 3329 4029 3341 4032
rect 3375 4029 3387 4063
rect 3329 4023 3387 4029
rect 3421 4063 3479 4069
rect 3421 4029 3433 4063
rect 3467 4060 3479 4063
rect 3878 4060 3884 4072
rect 3467 4032 3884 4060
rect 3467 4029 3479 4032
rect 3421 4023 3479 4029
rect 3878 4020 3884 4032
rect 3936 4020 3942 4072
rect 1104 3834 7544 3856
rect 1104 3782 2055 3834
rect 2107 3782 2119 3834
rect 2171 3782 2183 3834
rect 2235 3782 2247 3834
rect 2299 3782 4202 3834
rect 4254 3782 4266 3834
rect 4318 3782 4330 3834
rect 4382 3782 4394 3834
rect 4446 3782 6348 3834
rect 6400 3782 6412 3834
rect 6464 3782 6476 3834
rect 6528 3782 6540 3834
rect 6592 3782 7544 3834
rect 1104 3760 7544 3782
rect 3878 3720 3884 3732
rect 3839 3692 3884 3720
rect 3878 3680 3884 3692
rect 3936 3680 3942 3732
rect 5077 3723 5135 3729
rect 5077 3689 5089 3723
rect 5123 3720 5135 3723
rect 5626 3720 5632 3732
rect 5123 3692 5632 3720
rect 5123 3689 5135 3692
rect 5077 3683 5135 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 3786 3516 3792 3528
rect 3747 3488 3792 3516
rect 3786 3476 3792 3488
rect 3844 3476 3850 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5074 3516 5080 3528
rect 5031 3488 5080 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5074 3476 5080 3488
rect 5132 3476 5138 3528
rect 5166 3476 5172 3528
rect 5224 3525 5230 3528
rect 5224 3519 5237 3525
rect 5225 3516 5237 3519
rect 5810 3516 5816 3528
rect 5225 3488 5396 3516
rect 5771 3488 5816 3516
rect 5225 3485 5237 3488
rect 5224 3479 5237 3485
rect 5224 3476 5230 3479
rect 5368 3448 5396 3488
rect 5810 3476 5816 3488
rect 5868 3476 5874 3528
rect 5721 3451 5779 3457
rect 5721 3448 5733 3451
rect 5368 3420 5733 3448
rect 5721 3417 5733 3420
rect 5767 3417 5779 3451
rect 5721 3411 5779 3417
rect 1104 3290 7544 3312
rect 1104 3238 3128 3290
rect 3180 3238 3192 3290
rect 3244 3238 3256 3290
rect 3308 3238 3320 3290
rect 3372 3238 5275 3290
rect 5327 3238 5339 3290
rect 5391 3238 5403 3290
rect 5455 3238 5467 3290
rect 5519 3238 7544 3290
rect 1104 3216 7544 3238
rect 1104 2746 7544 2768
rect 1104 2694 2055 2746
rect 2107 2694 2119 2746
rect 2171 2694 2183 2746
rect 2235 2694 2247 2746
rect 2299 2694 4202 2746
rect 4254 2694 4266 2746
rect 4318 2694 4330 2746
rect 4382 2694 4394 2746
rect 4446 2694 6348 2746
rect 6400 2694 6412 2746
rect 6464 2694 6476 2746
rect 6528 2694 6540 2746
rect 6592 2694 7544 2746
rect 1104 2672 7544 2694
rect 1581 2635 1639 2641
rect 1581 2601 1593 2635
rect 1627 2632 1639 2635
rect 2774 2632 2780 2644
rect 1627 2604 2780 2632
rect 1627 2601 1639 2604
rect 1581 2595 1639 2601
rect 2774 2592 2780 2604
rect 2832 2592 2838 2644
rect 3237 2635 3295 2641
rect 3237 2601 3249 2635
rect 3283 2632 3295 2635
rect 3786 2632 3792 2644
rect 3283 2604 3792 2632
rect 3283 2601 3295 2604
rect 3237 2595 3295 2601
rect 3786 2592 3792 2604
rect 3844 2592 3850 2644
rect 4982 2592 4988 2644
rect 5040 2632 5046 2644
rect 5629 2635 5687 2641
rect 5629 2632 5641 2635
rect 5040 2604 5641 2632
rect 5040 2592 5046 2604
rect 5629 2601 5641 2604
rect 5675 2601 5687 2635
rect 5629 2595 5687 2601
rect 5810 2592 5816 2644
rect 5868 2632 5874 2644
rect 6641 2635 6699 2641
rect 6641 2632 6653 2635
rect 5868 2604 6653 2632
rect 5868 2592 5874 2604
rect 6641 2601 6653 2604
rect 6687 2601 6699 2635
rect 6641 2595 6699 2601
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 2958 2388 2964 2440
rect 3016 2428 3022 2440
rect 3053 2431 3111 2437
rect 3053 2428 3065 2431
rect 3016 2400 3065 2428
rect 3016 2388 3022 2400
rect 3053 2397 3065 2400
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 5813 2431 5871 2437
rect 5813 2397 5825 2431
rect 5859 2428 5871 2431
rect 5902 2428 5908 2440
rect 5859 2400 5908 2428
rect 5859 2397 5871 2400
rect 5813 2391 5871 2397
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 6822 2428 6828 2440
rect 6783 2400 6828 2428
rect 6822 2388 6828 2400
rect 6880 2388 6886 2440
rect 1104 2202 7544 2224
rect 1104 2150 3128 2202
rect 3180 2150 3192 2202
rect 3244 2150 3256 2202
rect 3308 2150 3320 2202
rect 3372 2150 5275 2202
rect 5327 2150 5339 2202
rect 5391 2150 5403 2202
rect 5455 2150 5467 2202
rect 5519 2150 7544 2202
rect 1104 2128 7544 2150
<< via1 >>
rect 2055 8134 2107 8186
rect 2119 8134 2171 8186
rect 2183 8134 2235 8186
rect 2247 8134 2299 8186
rect 4202 8134 4254 8186
rect 4266 8134 4318 8186
rect 4330 8134 4382 8186
rect 4394 8134 4446 8186
rect 6348 8134 6400 8186
rect 6412 8134 6464 8186
rect 6476 8134 6528 8186
rect 6540 8134 6592 8186
rect 4528 8032 4580 8084
rect 1308 7964 1360 8016
rect 4620 7828 4672 7880
rect 7196 7828 7248 7880
rect 4528 7803 4580 7812
rect 4528 7769 4537 7803
rect 4537 7769 4571 7803
rect 4571 7769 4580 7803
rect 4528 7760 4580 7769
rect 5632 7692 5684 7744
rect 3128 7590 3180 7642
rect 3192 7590 3244 7642
rect 3256 7590 3308 7642
rect 3320 7590 3372 7642
rect 5275 7590 5327 7642
rect 5339 7590 5391 7642
rect 5403 7590 5455 7642
rect 5467 7590 5519 7642
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 6828 7395 6880 7404
rect 6828 7361 6837 7395
rect 6837 7361 6871 7395
rect 6871 7361 6880 7395
rect 6828 7352 6880 7361
rect 4804 7148 4856 7200
rect 6644 7191 6696 7200
rect 6644 7157 6653 7191
rect 6653 7157 6687 7191
rect 6687 7157 6696 7191
rect 6644 7148 6696 7157
rect 2055 7046 2107 7098
rect 2119 7046 2171 7098
rect 2183 7046 2235 7098
rect 2247 7046 2299 7098
rect 4202 7046 4254 7098
rect 4266 7046 4318 7098
rect 4330 7046 4382 7098
rect 4394 7046 4446 7098
rect 6348 7046 6400 7098
rect 6412 7046 6464 7098
rect 6476 7046 6528 7098
rect 6540 7046 6592 7098
rect 3128 6502 3180 6554
rect 3192 6502 3244 6554
rect 3256 6502 3308 6554
rect 3320 6502 3372 6554
rect 5275 6502 5327 6554
rect 5339 6502 5391 6554
rect 5403 6502 5455 6554
rect 5467 6502 5519 6554
rect 2055 5958 2107 6010
rect 2119 5958 2171 6010
rect 2183 5958 2235 6010
rect 2247 5958 2299 6010
rect 4202 5958 4254 6010
rect 4266 5958 4318 6010
rect 4330 5958 4382 6010
rect 4394 5958 4446 6010
rect 6348 5958 6400 6010
rect 6412 5958 6464 6010
rect 6476 5958 6528 6010
rect 6540 5958 6592 6010
rect 4528 5856 4580 5908
rect 6644 5720 6696 5772
rect 4528 5652 4580 5704
rect 4620 5695 4672 5704
rect 4620 5661 4629 5695
rect 4629 5661 4663 5695
rect 4663 5661 4672 5695
rect 4620 5652 4672 5661
rect 4988 5652 5040 5704
rect 3424 5516 3476 5568
rect 5172 5516 5224 5568
rect 3128 5414 3180 5466
rect 3192 5414 3244 5466
rect 3256 5414 3308 5466
rect 3320 5414 3372 5466
rect 5275 5414 5327 5466
rect 5339 5414 5391 5466
rect 5403 5414 5455 5466
rect 5467 5414 5519 5466
rect 4528 5312 4580 5364
rect 3608 5219 3660 5228
rect 3056 5108 3108 5160
rect 3608 5185 3617 5219
rect 3617 5185 3651 5219
rect 3651 5185 3660 5219
rect 3608 5176 3660 5185
rect 3792 5176 3844 5228
rect 4896 5219 4948 5228
rect 4896 5185 4900 5219
rect 4900 5185 4934 5219
rect 4934 5185 4948 5219
rect 4896 5176 4948 5185
rect 4068 4972 4120 5024
rect 4528 4972 4580 5024
rect 5448 5176 5500 5228
rect 4988 5040 5040 5092
rect 5632 4972 5684 5024
rect 2055 4870 2107 4922
rect 2119 4870 2171 4922
rect 2183 4870 2235 4922
rect 2247 4870 2299 4922
rect 4202 4870 4254 4922
rect 4266 4870 4318 4922
rect 4330 4870 4382 4922
rect 4394 4870 4446 4922
rect 6348 4870 6400 4922
rect 6412 4870 6464 4922
rect 6476 4870 6528 4922
rect 6540 4870 6592 4922
rect 4528 4768 4580 4820
rect 4896 4811 4948 4820
rect 4896 4777 4905 4811
rect 4905 4777 4939 4811
rect 4939 4777 4948 4811
rect 4896 4768 4948 4777
rect 2964 4632 3016 4684
rect 1400 4607 1452 4616
rect 1400 4573 1409 4607
rect 1409 4573 1443 4607
rect 1443 4573 1452 4607
rect 1400 4564 1452 4573
rect 3608 4564 3660 4616
rect 3884 4564 3936 4616
rect 4068 4607 4120 4616
rect 4068 4573 4077 4607
rect 4077 4573 4111 4607
rect 4111 4573 4120 4607
rect 4344 4607 4396 4616
rect 4068 4564 4120 4573
rect 4344 4573 4353 4607
rect 4353 4573 4387 4607
rect 4387 4573 4396 4607
rect 4344 4564 4396 4573
rect 4804 4700 4856 4752
rect 5448 4700 5500 4752
rect 5172 4632 5224 4684
rect 5080 4607 5132 4616
rect 5080 4573 5089 4607
rect 5089 4573 5123 4607
rect 5123 4573 5132 4607
rect 5080 4564 5132 4573
rect 5632 4607 5684 4616
rect 2780 4539 2832 4548
rect 2780 4505 2789 4539
rect 2789 4505 2823 4539
rect 2823 4505 2832 4539
rect 2780 4496 2832 4505
rect 3056 4539 3108 4548
rect 3056 4505 3065 4539
rect 3065 4505 3099 4539
rect 3099 4505 3108 4539
rect 3056 4496 3108 4505
rect 3516 4496 3568 4548
rect 5172 4496 5224 4548
rect 5632 4573 5641 4607
rect 5641 4573 5675 4607
rect 5675 4573 5684 4607
rect 5632 4564 5684 4573
rect 3424 4428 3476 4480
rect 4620 4428 4672 4480
rect 6736 4471 6788 4480
rect 6736 4437 6745 4471
rect 6745 4437 6779 4471
rect 6779 4437 6788 4471
rect 6736 4428 6788 4437
rect 3128 4326 3180 4378
rect 3192 4326 3244 4378
rect 3256 4326 3308 4378
rect 3320 4326 3372 4378
rect 5275 4326 5327 4378
rect 5339 4326 5391 4378
rect 5403 4326 5455 4378
rect 5467 4326 5519 4378
rect 3792 4267 3844 4276
rect 3792 4233 3801 4267
rect 3801 4233 3835 4267
rect 3835 4233 3844 4267
rect 3792 4224 3844 4233
rect 4344 4224 4396 4276
rect 2964 4088 3016 4140
rect 3424 4156 3476 4208
rect 5080 4156 5132 4208
rect 3516 4088 3568 4140
rect 4896 4131 4948 4140
rect 4896 4097 4905 4131
rect 4905 4097 4939 4131
rect 4939 4097 4948 4131
rect 4896 4088 4948 4097
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 2780 4020 2832 4072
rect 3884 4020 3936 4072
rect 2055 3782 2107 3834
rect 2119 3782 2171 3834
rect 2183 3782 2235 3834
rect 2247 3782 2299 3834
rect 4202 3782 4254 3834
rect 4266 3782 4318 3834
rect 4330 3782 4382 3834
rect 4394 3782 4446 3834
rect 6348 3782 6400 3834
rect 6412 3782 6464 3834
rect 6476 3782 6528 3834
rect 6540 3782 6592 3834
rect 3884 3723 3936 3732
rect 3884 3689 3893 3723
rect 3893 3689 3927 3723
rect 3927 3689 3936 3723
rect 3884 3680 3936 3689
rect 5632 3680 5684 3732
rect 3792 3519 3844 3528
rect 3792 3485 3801 3519
rect 3801 3485 3835 3519
rect 3835 3485 3844 3519
rect 3792 3476 3844 3485
rect 5080 3476 5132 3528
rect 5172 3519 5224 3528
rect 5172 3485 5191 3519
rect 5191 3485 5224 3519
rect 5816 3519 5868 3528
rect 5172 3476 5224 3485
rect 5816 3485 5825 3519
rect 5825 3485 5859 3519
rect 5859 3485 5868 3519
rect 5816 3476 5868 3485
rect 3128 3238 3180 3290
rect 3192 3238 3244 3290
rect 3256 3238 3308 3290
rect 3320 3238 3372 3290
rect 5275 3238 5327 3290
rect 5339 3238 5391 3290
rect 5403 3238 5455 3290
rect 5467 3238 5519 3290
rect 2055 2694 2107 2746
rect 2119 2694 2171 2746
rect 2183 2694 2235 2746
rect 2247 2694 2299 2746
rect 4202 2694 4254 2746
rect 4266 2694 4318 2746
rect 4330 2694 4382 2746
rect 4394 2694 4446 2746
rect 6348 2694 6400 2746
rect 6412 2694 6464 2746
rect 6476 2694 6528 2746
rect 6540 2694 6592 2746
rect 2780 2592 2832 2644
rect 3792 2592 3844 2644
rect 4988 2592 5040 2644
rect 5816 2592 5868 2644
rect 20 2388 72 2440
rect 2964 2388 3016 2440
rect 5908 2388 5960 2440
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 3128 2150 3180 2202
rect 3192 2150 3244 2202
rect 3256 2150 3308 2202
rect 3320 2150 3372 2202
rect 5275 2150 5327 2202
rect 5339 2150 5391 2202
rect 5403 2150 5455 2202
rect 5467 2150 5519 2202
<< metal2 >>
rect 1306 10074 1362 10874
rect 4250 10074 4306 10874
rect 4356 10118 4568 10146
rect 1320 8022 1348 10074
rect 4264 10010 4292 10074
rect 4356 10010 4384 10118
rect 4264 9982 4384 10010
rect 1398 8528 1454 8537
rect 1398 8463 1454 8472
rect 1308 8016 1360 8022
rect 1308 7958 1360 7964
rect 1412 7410 1440 8463
rect 2029 8188 2325 8208
rect 2085 8186 2109 8188
rect 2165 8186 2189 8188
rect 2245 8186 2269 8188
rect 2107 8134 2109 8186
rect 2171 8134 2183 8186
rect 2245 8134 2247 8186
rect 2085 8132 2109 8134
rect 2165 8132 2189 8134
rect 2245 8132 2269 8134
rect 2029 8112 2325 8132
rect 4176 8188 4472 8208
rect 4232 8186 4256 8188
rect 4312 8186 4336 8188
rect 4392 8186 4416 8188
rect 4254 8134 4256 8186
rect 4318 8134 4330 8186
rect 4392 8134 4394 8186
rect 4232 8132 4256 8134
rect 4312 8132 4336 8134
rect 4392 8132 4416 8134
rect 4176 8112 4472 8132
rect 4540 8090 4568 10118
rect 7194 10074 7250 10874
rect 6826 8800 6882 8809
rect 6826 8735 6882 8744
rect 6322 8188 6618 8208
rect 6378 8186 6402 8188
rect 6458 8186 6482 8188
rect 6538 8186 6562 8188
rect 6400 8134 6402 8186
rect 6464 8134 6476 8186
rect 6538 8134 6540 8186
rect 6378 8132 6402 8134
rect 6458 8132 6482 8134
rect 6538 8132 6562 8134
rect 6322 8112 6618 8132
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4620 7880 4672 7886
rect 4620 7822 4672 7828
rect 4528 7812 4580 7818
rect 4528 7754 4580 7760
rect 3102 7644 3398 7664
rect 3158 7642 3182 7644
rect 3238 7642 3262 7644
rect 3318 7642 3342 7644
rect 3180 7590 3182 7642
rect 3244 7590 3256 7642
rect 3318 7590 3320 7642
rect 3158 7588 3182 7590
rect 3238 7588 3262 7590
rect 3318 7588 3342 7590
rect 3102 7568 3398 7588
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 2029 7100 2325 7120
rect 2085 7098 2109 7100
rect 2165 7098 2189 7100
rect 2245 7098 2269 7100
rect 2107 7046 2109 7098
rect 2171 7046 2183 7098
rect 2245 7046 2247 7098
rect 2085 7044 2109 7046
rect 2165 7044 2189 7046
rect 2245 7044 2269 7046
rect 2029 7024 2325 7044
rect 4176 7100 4472 7120
rect 4232 7098 4256 7100
rect 4312 7098 4336 7100
rect 4392 7098 4416 7100
rect 4254 7046 4256 7098
rect 4318 7046 4330 7098
rect 4392 7046 4394 7098
rect 4232 7044 4256 7046
rect 4312 7044 4336 7046
rect 4392 7044 4416 7046
rect 4176 7024 4472 7044
rect 3102 6556 3398 6576
rect 3158 6554 3182 6556
rect 3238 6554 3262 6556
rect 3318 6554 3342 6556
rect 3180 6502 3182 6554
rect 3244 6502 3256 6554
rect 3318 6502 3320 6554
rect 3158 6500 3182 6502
rect 3238 6500 3262 6502
rect 3318 6500 3342 6502
rect 3102 6480 3398 6500
rect 2029 6012 2325 6032
rect 2085 6010 2109 6012
rect 2165 6010 2189 6012
rect 2245 6010 2269 6012
rect 2107 5958 2109 6010
rect 2171 5958 2183 6010
rect 2245 5958 2247 6010
rect 2085 5956 2109 5958
rect 2165 5956 2189 5958
rect 2245 5956 2269 5958
rect 2029 5936 2325 5956
rect 4176 6012 4472 6032
rect 4232 6010 4256 6012
rect 4312 6010 4336 6012
rect 4392 6010 4416 6012
rect 4254 5958 4256 6010
rect 4318 5958 4330 6010
rect 4392 5958 4394 6010
rect 4232 5956 4256 5958
rect 4312 5956 4336 5958
rect 4392 5956 4416 5958
rect 4176 5936 4472 5956
rect 4540 5914 4568 7754
rect 4528 5908 4580 5914
rect 4528 5850 4580 5856
rect 4632 5794 4660 7822
rect 5632 7744 5684 7750
rect 5632 7686 5684 7692
rect 5249 7644 5545 7664
rect 5305 7642 5329 7644
rect 5385 7642 5409 7644
rect 5465 7642 5489 7644
rect 5327 7590 5329 7642
rect 5391 7590 5403 7642
rect 5465 7590 5467 7642
rect 5305 7588 5329 7590
rect 5385 7588 5409 7590
rect 5465 7588 5489 7590
rect 5249 7568 5545 7588
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4540 5766 4660 5794
rect 4540 5710 4568 5766
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4620 5704 4672 5710
rect 4620 5646 4672 5652
rect 3424 5568 3476 5574
rect 3424 5510 3476 5516
rect 3102 5468 3398 5488
rect 3158 5466 3182 5468
rect 3238 5466 3262 5468
rect 3318 5466 3342 5468
rect 3180 5414 3182 5466
rect 3244 5414 3256 5466
rect 3318 5414 3320 5466
rect 3158 5412 3182 5414
rect 3238 5412 3262 5414
rect 3318 5412 3342 5414
rect 3102 5392 3398 5412
rect 3056 5160 3108 5166
rect 3056 5102 3108 5108
rect 2029 4924 2325 4944
rect 2085 4922 2109 4924
rect 2165 4922 2189 4924
rect 2245 4922 2269 4924
rect 2107 4870 2109 4922
rect 2171 4870 2183 4922
rect 2245 4870 2247 4922
rect 2085 4868 2109 4870
rect 2165 4868 2189 4870
rect 2245 4868 2269 4870
rect 2029 4848 2325 4868
rect 2964 4684 3016 4690
rect 2964 4626 3016 4632
rect 1400 4616 1452 4622
rect 1400 4558 1452 4564
rect 1412 4185 1440 4558
rect 2780 4548 2832 4554
rect 2780 4490 2832 4496
rect 1398 4176 1454 4185
rect 1398 4111 1454 4120
rect 2792 4078 2820 4490
rect 2976 4146 3004 4626
rect 3068 4554 3096 5102
rect 3056 4548 3108 4554
rect 3056 4490 3108 4496
rect 3436 4486 3464 5510
rect 4540 5370 4568 5646
rect 4528 5364 4580 5370
rect 4528 5306 4580 5312
rect 3608 5228 3660 5234
rect 3608 5170 3660 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3620 4622 3648 5170
rect 3608 4616 3660 4622
rect 3608 4558 3660 4564
rect 3516 4548 3568 4554
rect 3516 4490 3568 4496
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3102 4380 3398 4400
rect 3158 4378 3182 4380
rect 3238 4378 3262 4380
rect 3318 4378 3342 4380
rect 3180 4326 3182 4378
rect 3244 4326 3256 4378
rect 3318 4326 3320 4378
rect 3158 4324 3182 4326
rect 3238 4324 3262 4326
rect 3318 4324 3342 4326
rect 3102 4304 3398 4324
rect 3436 4214 3464 4422
rect 3424 4208 3476 4214
rect 3424 4150 3476 4156
rect 3528 4146 3556 4490
rect 3804 4282 3832 5170
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4080 4622 4108 4966
rect 4176 4924 4472 4944
rect 4232 4922 4256 4924
rect 4312 4922 4336 4924
rect 4392 4922 4416 4924
rect 4254 4870 4256 4922
rect 4318 4870 4330 4922
rect 4392 4870 4394 4922
rect 4232 4868 4256 4870
rect 4312 4868 4336 4870
rect 4392 4868 4416 4870
rect 4176 4848 4472 4868
rect 4540 4826 4568 4966
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 4068 4616 4120 4622
rect 4068 4558 4120 4564
rect 4344 4616 4396 4622
rect 4344 4558 4396 4564
rect 3792 4276 3844 4282
rect 3792 4218 3844 4224
rect 2964 4140 3016 4146
rect 2964 4082 3016 4088
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3896 4078 3924 4558
rect 4356 4282 4384 4558
rect 4632 4486 4660 5646
rect 4816 4758 4844 7142
rect 5249 6556 5545 6576
rect 5305 6554 5329 6556
rect 5385 6554 5409 6556
rect 5465 6554 5489 6556
rect 5327 6502 5329 6554
rect 5391 6502 5403 6554
rect 5465 6502 5467 6554
rect 5305 6500 5329 6502
rect 5385 6500 5409 6502
rect 5465 6500 5489 6502
rect 5249 6480 5545 6500
rect 4988 5704 5040 5710
rect 4988 5646 5040 5652
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4908 4826 4936 5170
rect 5000 5098 5028 5646
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4988 5092 5040 5098
rect 4988 5034 5040 5040
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 4620 4480 4672 4486
rect 4620 4422 4672 4428
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 4908 4146 4936 4762
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 3884 4072 3936 4078
rect 3884 4014 3936 4020
rect 2029 3836 2325 3856
rect 2085 3834 2109 3836
rect 2165 3834 2189 3836
rect 2245 3834 2269 3836
rect 2107 3782 2109 3834
rect 2171 3782 2183 3834
rect 2245 3782 2247 3834
rect 2085 3780 2109 3782
rect 2165 3780 2189 3782
rect 2245 3780 2269 3782
rect 2029 3760 2325 3780
rect 2029 2748 2325 2768
rect 2085 2746 2109 2748
rect 2165 2746 2189 2748
rect 2245 2746 2269 2748
rect 2107 2694 2109 2746
rect 2171 2694 2183 2746
rect 2245 2694 2247 2746
rect 2085 2692 2109 2694
rect 2165 2692 2189 2694
rect 2245 2692 2269 2694
rect 2029 2672 2325 2692
rect 2792 2650 2820 4014
rect 3896 3738 3924 4014
rect 4176 3836 4472 3856
rect 4232 3834 4256 3836
rect 4312 3834 4336 3836
rect 4392 3834 4416 3836
rect 4254 3782 4256 3834
rect 4318 3782 4330 3834
rect 4392 3782 4394 3834
rect 4232 3780 4256 3782
rect 4312 3780 4336 3782
rect 4392 3780 4416 3782
rect 4176 3760 4472 3780
rect 3884 3732 3936 3738
rect 3884 3674 3936 3680
rect 3792 3528 3844 3534
rect 3792 3470 3844 3476
rect 3102 3292 3398 3312
rect 3158 3290 3182 3292
rect 3238 3290 3262 3292
rect 3318 3290 3342 3292
rect 3180 3238 3182 3290
rect 3244 3238 3256 3290
rect 3318 3238 3320 3290
rect 3158 3236 3182 3238
rect 3238 3236 3262 3238
rect 3318 3236 3342 3238
rect 3102 3216 3398 3236
rect 3804 2650 3832 3470
rect 4176 2748 4472 2768
rect 4232 2746 4256 2748
rect 4312 2746 4336 2748
rect 4392 2746 4416 2748
rect 4254 2694 4256 2746
rect 4318 2694 4330 2746
rect 4392 2694 4394 2746
rect 4232 2692 4256 2694
rect 4312 2692 4336 2694
rect 4392 2692 4416 2694
rect 4176 2672 4472 2692
rect 5000 2650 5028 5034
rect 5184 4690 5212 5510
rect 5249 5468 5545 5488
rect 5305 5466 5329 5468
rect 5385 5466 5409 5468
rect 5465 5466 5489 5468
rect 5327 5414 5329 5466
rect 5391 5414 5403 5466
rect 5465 5414 5467 5466
rect 5305 5412 5329 5414
rect 5385 5412 5409 5414
rect 5465 5412 5489 5414
rect 5249 5392 5545 5412
rect 5448 5228 5500 5234
rect 5448 5170 5500 5176
rect 5460 4758 5488 5170
rect 5644 5030 5672 7686
rect 6840 7410 6868 8735
rect 7208 7886 7236 10074
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 6644 7200 6696 7206
rect 6644 7142 6696 7148
rect 6322 7100 6618 7120
rect 6378 7098 6402 7100
rect 6458 7098 6482 7100
rect 6538 7098 6562 7100
rect 6400 7046 6402 7098
rect 6464 7046 6476 7098
rect 6538 7046 6540 7098
rect 6378 7044 6402 7046
rect 6458 7044 6482 7046
rect 6538 7044 6562 7046
rect 6322 7024 6618 7044
rect 6322 6012 6618 6032
rect 6378 6010 6402 6012
rect 6458 6010 6482 6012
rect 6538 6010 6562 6012
rect 6400 5958 6402 6010
rect 6464 5958 6476 6010
rect 6538 5958 6540 6010
rect 6378 5956 6402 5958
rect 6458 5956 6482 5958
rect 6538 5956 6562 5958
rect 6322 5936 6618 5956
rect 6656 5778 6684 7142
rect 6644 5772 6696 5778
rect 6644 5714 6696 5720
rect 5632 5024 5684 5030
rect 5632 4966 5684 4972
rect 6322 4924 6618 4944
rect 6378 4922 6402 4924
rect 6458 4922 6482 4924
rect 6538 4922 6562 4924
rect 6400 4870 6402 4922
rect 6464 4870 6476 4922
rect 6538 4870 6540 4922
rect 6378 4868 6402 4870
rect 6458 4868 6482 4870
rect 6538 4868 6562 4870
rect 6322 4848 6618 4868
rect 5448 4752 5500 4758
rect 5448 4694 5500 4700
rect 5172 4684 5224 4690
rect 5172 4626 5224 4632
rect 5080 4616 5132 4622
rect 5080 4558 5132 4564
rect 5632 4616 5684 4622
rect 5632 4558 5684 4564
rect 5092 4214 5120 4558
rect 5172 4548 5224 4554
rect 5172 4490 5224 4496
rect 5080 4208 5132 4214
rect 5080 4150 5132 4156
rect 5092 3534 5120 4150
rect 5184 4146 5212 4490
rect 5249 4380 5545 4400
rect 5305 4378 5329 4380
rect 5385 4378 5409 4380
rect 5465 4378 5489 4380
rect 5327 4326 5329 4378
rect 5391 4326 5403 4378
rect 5465 4326 5467 4378
rect 5305 4324 5329 4326
rect 5385 4324 5409 4326
rect 5465 4324 5489 4326
rect 5249 4304 5545 4324
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5184 3534 5212 4082
rect 5644 3738 5672 4558
rect 6736 4480 6788 4486
rect 6734 4448 6736 4457
rect 6788 4448 6790 4457
rect 6734 4383 6790 4392
rect 6322 3836 6618 3856
rect 6378 3834 6402 3836
rect 6458 3834 6482 3836
rect 6538 3834 6562 3836
rect 6400 3782 6402 3834
rect 6464 3782 6476 3834
rect 6538 3782 6540 3834
rect 6378 3780 6402 3782
rect 6458 3780 6482 3782
rect 6538 3780 6562 3782
rect 6322 3760 6618 3780
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5080 3528 5132 3534
rect 5080 3470 5132 3476
rect 5172 3528 5224 3534
rect 5172 3470 5224 3476
rect 5816 3528 5868 3534
rect 5816 3470 5868 3476
rect 5249 3292 5545 3312
rect 5305 3290 5329 3292
rect 5385 3290 5409 3292
rect 5465 3290 5489 3292
rect 5327 3238 5329 3290
rect 5391 3238 5403 3290
rect 5465 3238 5467 3290
rect 5305 3236 5329 3238
rect 5385 3236 5409 3238
rect 5465 3236 5489 3238
rect 5249 3216 5545 3236
rect 5828 2650 5856 3470
rect 6322 2748 6618 2768
rect 6378 2746 6402 2748
rect 6458 2746 6482 2748
rect 6538 2746 6562 2748
rect 6400 2694 6402 2746
rect 6464 2694 6476 2746
rect 6538 2694 6540 2746
rect 6378 2692 6402 2694
rect 6458 2692 6482 2694
rect 6538 2692 6562 2694
rect 6322 2672 6618 2692
rect 2780 2644 2832 2650
rect 2780 2586 2832 2592
rect 3792 2644 3844 2650
rect 3792 2586 3844 2592
rect 4988 2644 5040 2650
rect 4988 2586 5040 2592
rect 5816 2644 5868 2650
rect 5816 2586 5868 2592
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 5908 2440 5960 2446
rect 5908 2382 5960 2388
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 32 800 60 2382
rect 2976 800 3004 2382
rect 3102 2204 3398 2224
rect 3158 2202 3182 2204
rect 3238 2202 3262 2204
rect 3318 2202 3342 2204
rect 3180 2150 3182 2202
rect 3244 2150 3256 2202
rect 3318 2150 3320 2202
rect 3158 2148 3182 2150
rect 3238 2148 3262 2150
rect 3318 2148 3342 2150
rect 3102 2128 3398 2148
rect 5249 2204 5545 2224
rect 5305 2202 5329 2204
rect 5385 2202 5409 2204
rect 5465 2202 5489 2204
rect 5327 2150 5329 2202
rect 5391 2150 5403 2202
rect 5465 2150 5467 2202
rect 5305 2148 5329 2150
rect 5385 2148 5409 2150
rect 5465 2148 5489 2150
rect 5249 2128 5545 2148
rect 5920 800 5948 2382
rect 18 0 74 800
rect 2962 0 3018 800
rect 5906 0 5962 800
rect 6840 105 6868 2382
rect 6826 96 6882 105
rect 6826 31 6882 40
<< via2 >>
rect 1398 8472 1454 8528
rect 2029 8186 2085 8188
rect 2109 8186 2165 8188
rect 2189 8186 2245 8188
rect 2269 8186 2325 8188
rect 2029 8134 2055 8186
rect 2055 8134 2085 8186
rect 2109 8134 2119 8186
rect 2119 8134 2165 8186
rect 2189 8134 2235 8186
rect 2235 8134 2245 8186
rect 2269 8134 2299 8186
rect 2299 8134 2325 8186
rect 2029 8132 2085 8134
rect 2109 8132 2165 8134
rect 2189 8132 2245 8134
rect 2269 8132 2325 8134
rect 4176 8186 4232 8188
rect 4256 8186 4312 8188
rect 4336 8186 4392 8188
rect 4416 8186 4472 8188
rect 4176 8134 4202 8186
rect 4202 8134 4232 8186
rect 4256 8134 4266 8186
rect 4266 8134 4312 8186
rect 4336 8134 4382 8186
rect 4382 8134 4392 8186
rect 4416 8134 4446 8186
rect 4446 8134 4472 8186
rect 4176 8132 4232 8134
rect 4256 8132 4312 8134
rect 4336 8132 4392 8134
rect 4416 8132 4472 8134
rect 6826 8744 6882 8800
rect 6322 8186 6378 8188
rect 6402 8186 6458 8188
rect 6482 8186 6538 8188
rect 6562 8186 6618 8188
rect 6322 8134 6348 8186
rect 6348 8134 6378 8186
rect 6402 8134 6412 8186
rect 6412 8134 6458 8186
rect 6482 8134 6528 8186
rect 6528 8134 6538 8186
rect 6562 8134 6592 8186
rect 6592 8134 6618 8186
rect 6322 8132 6378 8134
rect 6402 8132 6458 8134
rect 6482 8132 6538 8134
rect 6562 8132 6618 8134
rect 3102 7642 3158 7644
rect 3182 7642 3238 7644
rect 3262 7642 3318 7644
rect 3342 7642 3398 7644
rect 3102 7590 3128 7642
rect 3128 7590 3158 7642
rect 3182 7590 3192 7642
rect 3192 7590 3238 7642
rect 3262 7590 3308 7642
rect 3308 7590 3318 7642
rect 3342 7590 3372 7642
rect 3372 7590 3398 7642
rect 3102 7588 3158 7590
rect 3182 7588 3238 7590
rect 3262 7588 3318 7590
rect 3342 7588 3398 7590
rect 2029 7098 2085 7100
rect 2109 7098 2165 7100
rect 2189 7098 2245 7100
rect 2269 7098 2325 7100
rect 2029 7046 2055 7098
rect 2055 7046 2085 7098
rect 2109 7046 2119 7098
rect 2119 7046 2165 7098
rect 2189 7046 2235 7098
rect 2235 7046 2245 7098
rect 2269 7046 2299 7098
rect 2299 7046 2325 7098
rect 2029 7044 2085 7046
rect 2109 7044 2165 7046
rect 2189 7044 2245 7046
rect 2269 7044 2325 7046
rect 4176 7098 4232 7100
rect 4256 7098 4312 7100
rect 4336 7098 4392 7100
rect 4416 7098 4472 7100
rect 4176 7046 4202 7098
rect 4202 7046 4232 7098
rect 4256 7046 4266 7098
rect 4266 7046 4312 7098
rect 4336 7046 4382 7098
rect 4382 7046 4392 7098
rect 4416 7046 4446 7098
rect 4446 7046 4472 7098
rect 4176 7044 4232 7046
rect 4256 7044 4312 7046
rect 4336 7044 4392 7046
rect 4416 7044 4472 7046
rect 3102 6554 3158 6556
rect 3182 6554 3238 6556
rect 3262 6554 3318 6556
rect 3342 6554 3398 6556
rect 3102 6502 3128 6554
rect 3128 6502 3158 6554
rect 3182 6502 3192 6554
rect 3192 6502 3238 6554
rect 3262 6502 3308 6554
rect 3308 6502 3318 6554
rect 3342 6502 3372 6554
rect 3372 6502 3398 6554
rect 3102 6500 3158 6502
rect 3182 6500 3238 6502
rect 3262 6500 3318 6502
rect 3342 6500 3398 6502
rect 2029 6010 2085 6012
rect 2109 6010 2165 6012
rect 2189 6010 2245 6012
rect 2269 6010 2325 6012
rect 2029 5958 2055 6010
rect 2055 5958 2085 6010
rect 2109 5958 2119 6010
rect 2119 5958 2165 6010
rect 2189 5958 2235 6010
rect 2235 5958 2245 6010
rect 2269 5958 2299 6010
rect 2299 5958 2325 6010
rect 2029 5956 2085 5958
rect 2109 5956 2165 5958
rect 2189 5956 2245 5958
rect 2269 5956 2325 5958
rect 4176 6010 4232 6012
rect 4256 6010 4312 6012
rect 4336 6010 4392 6012
rect 4416 6010 4472 6012
rect 4176 5958 4202 6010
rect 4202 5958 4232 6010
rect 4256 5958 4266 6010
rect 4266 5958 4312 6010
rect 4336 5958 4382 6010
rect 4382 5958 4392 6010
rect 4416 5958 4446 6010
rect 4446 5958 4472 6010
rect 4176 5956 4232 5958
rect 4256 5956 4312 5958
rect 4336 5956 4392 5958
rect 4416 5956 4472 5958
rect 5249 7642 5305 7644
rect 5329 7642 5385 7644
rect 5409 7642 5465 7644
rect 5489 7642 5545 7644
rect 5249 7590 5275 7642
rect 5275 7590 5305 7642
rect 5329 7590 5339 7642
rect 5339 7590 5385 7642
rect 5409 7590 5455 7642
rect 5455 7590 5465 7642
rect 5489 7590 5519 7642
rect 5519 7590 5545 7642
rect 5249 7588 5305 7590
rect 5329 7588 5385 7590
rect 5409 7588 5465 7590
rect 5489 7588 5545 7590
rect 3102 5466 3158 5468
rect 3182 5466 3238 5468
rect 3262 5466 3318 5468
rect 3342 5466 3398 5468
rect 3102 5414 3128 5466
rect 3128 5414 3158 5466
rect 3182 5414 3192 5466
rect 3192 5414 3238 5466
rect 3262 5414 3308 5466
rect 3308 5414 3318 5466
rect 3342 5414 3372 5466
rect 3372 5414 3398 5466
rect 3102 5412 3158 5414
rect 3182 5412 3238 5414
rect 3262 5412 3318 5414
rect 3342 5412 3398 5414
rect 2029 4922 2085 4924
rect 2109 4922 2165 4924
rect 2189 4922 2245 4924
rect 2269 4922 2325 4924
rect 2029 4870 2055 4922
rect 2055 4870 2085 4922
rect 2109 4870 2119 4922
rect 2119 4870 2165 4922
rect 2189 4870 2235 4922
rect 2235 4870 2245 4922
rect 2269 4870 2299 4922
rect 2299 4870 2325 4922
rect 2029 4868 2085 4870
rect 2109 4868 2165 4870
rect 2189 4868 2245 4870
rect 2269 4868 2325 4870
rect 1398 4120 1454 4176
rect 3102 4378 3158 4380
rect 3182 4378 3238 4380
rect 3262 4378 3318 4380
rect 3342 4378 3398 4380
rect 3102 4326 3128 4378
rect 3128 4326 3158 4378
rect 3182 4326 3192 4378
rect 3192 4326 3238 4378
rect 3262 4326 3308 4378
rect 3308 4326 3318 4378
rect 3342 4326 3372 4378
rect 3372 4326 3398 4378
rect 3102 4324 3158 4326
rect 3182 4324 3238 4326
rect 3262 4324 3318 4326
rect 3342 4324 3398 4326
rect 4176 4922 4232 4924
rect 4256 4922 4312 4924
rect 4336 4922 4392 4924
rect 4416 4922 4472 4924
rect 4176 4870 4202 4922
rect 4202 4870 4232 4922
rect 4256 4870 4266 4922
rect 4266 4870 4312 4922
rect 4336 4870 4382 4922
rect 4382 4870 4392 4922
rect 4416 4870 4446 4922
rect 4446 4870 4472 4922
rect 4176 4868 4232 4870
rect 4256 4868 4312 4870
rect 4336 4868 4392 4870
rect 4416 4868 4472 4870
rect 5249 6554 5305 6556
rect 5329 6554 5385 6556
rect 5409 6554 5465 6556
rect 5489 6554 5545 6556
rect 5249 6502 5275 6554
rect 5275 6502 5305 6554
rect 5329 6502 5339 6554
rect 5339 6502 5385 6554
rect 5409 6502 5455 6554
rect 5455 6502 5465 6554
rect 5489 6502 5519 6554
rect 5519 6502 5545 6554
rect 5249 6500 5305 6502
rect 5329 6500 5385 6502
rect 5409 6500 5465 6502
rect 5489 6500 5545 6502
rect 2029 3834 2085 3836
rect 2109 3834 2165 3836
rect 2189 3834 2245 3836
rect 2269 3834 2325 3836
rect 2029 3782 2055 3834
rect 2055 3782 2085 3834
rect 2109 3782 2119 3834
rect 2119 3782 2165 3834
rect 2189 3782 2235 3834
rect 2235 3782 2245 3834
rect 2269 3782 2299 3834
rect 2299 3782 2325 3834
rect 2029 3780 2085 3782
rect 2109 3780 2165 3782
rect 2189 3780 2245 3782
rect 2269 3780 2325 3782
rect 2029 2746 2085 2748
rect 2109 2746 2165 2748
rect 2189 2746 2245 2748
rect 2269 2746 2325 2748
rect 2029 2694 2055 2746
rect 2055 2694 2085 2746
rect 2109 2694 2119 2746
rect 2119 2694 2165 2746
rect 2189 2694 2235 2746
rect 2235 2694 2245 2746
rect 2269 2694 2299 2746
rect 2299 2694 2325 2746
rect 2029 2692 2085 2694
rect 2109 2692 2165 2694
rect 2189 2692 2245 2694
rect 2269 2692 2325 2694
rect 4176 3834 4232 3836
rect 4256 3834 4312 3836
rect 4336 3834 4392 3836
rect 4416 3834 4472 3836
rect 4176 3782 4202 3834
rect 4202 3782 4232 3834
rect 4256 3782 4266 3834
rect 4266 3782 4312 3834
rect 4336 3782 4382 3834
rect 4382 3782 4392 3834
rect 4416 3782 4446 3834
rect 4446 3782 4472 3834
rect 4176 3780 4232 3782
rect 4256 3780 4312 3782
rect 4336 3780 4392 3782
rect 4416 3780 4472 3782
rect 3102 3290 3158 3292
rect 3182 3290 3238 3292
rect 3262 3290 3318 3292
rect 3342 3290 3398 3292
rect 3102 3238 3128 3290
rect 3128 3238 3158 3290
rect 3182 3238 3192 3290
rect 3192 3238 3238 3290
rect 3262 3238 3308 3290
rect 3308 3238 3318 3290
rect 3342 3238 3372 3290
rect 3372 3238 3398 3290
rect 3102 3236 3158 3238
rect 3182 3236 3238 3238
rect 3262 3236 3318 3238
rect 3342 3236 3398 3238
rect 4176 2746 4232 2748
rect 4256 2746 4312 2748
rect 4336 2746 4392 2748
rect 4416 2746 4472 2748
rect 4176 2694 4202 2746
rect 4202 2694 4232 2746
rect 4256 2694 4266 2746
rect 4266 2694 4312 2746
rect 4336 2694 4382 2746
rect 4382 2694 4392 2746
rect 4416 2694 4446 2746
rect 4446 2694 4472 2746
rect 4176 2692 4232 2694
rect 4256 2692 4312 2694
rect 4336 2692 4392 2694
rect 4416 2692 4472 2694
rect 5249 5466 5305 5468
rect 5329 5466 5385 5468
rect 5409 5466 5465 5468
rect 5489 5466 5545 5468
rect 5249 5414 5275 5466
rect 5275 5414 5305 5466
rect 5329 5414 5339 5466
rect 5339 5414 5385 5466
rect 5409 5414 5455 5466
rect 5455 5414 5465 5466
rect 5489 5414 5519 5466
rect 5519 5414 5545 5466
rect 5249 5412 5305 5414
rect 5329 5412 5385 5414
rect 5409 5412 5465 5414
rect 5489 5412 5545 5414
rect 6322 7098 6378 7100
rect 6402 7098 6458 7100
rect 6482 7098 6538 7100
rect 6562 7098 6618 7100
rect 6322 7046 6348 7098
rect 6348 7046 6378 7098
rect 6402 7046 6412 7098
rect 6412 7046 6458 7098
rect 6482 7046 6528 7098
rect 6528 7046 6538 7098
rect 6562 7046 6592 7098
rect 6592 7046 6618 7098
rect 6322 7044 6378 7046
rect 6402 7044 6458 7046
rect 6482 7044 6538 7046
rect 6562 7044 6618 7046
rect 6322 6010 6378 6012
rect 6402 6010 6458 6012
rect 6482 6010 6538 6012
rect 6562 6010 6618 6012
rect 6322 5958 6348 6010
rect 6348 5958 6378 6010
rect 6402 5958 6412 6010
rect 6412 5958 6458 6010
rect 6482 5958 6528 6010
rect 6528 5958 6538 6010
rect 6562 5958 6592 6010
rect 6592 5958 6618 6010
rect 6322 5956 6378 5958
rect 6402 5956 6458 5958
rect 6482 5956 6538 5958
rect 6562 5956 6618 5958
rect 6322 4922 6378 4924
rect 6402 4922 6458 4924
rect 6482 4922 6538 4924
rect 6562 4922 6618 4924
rect 6322 4870 6348 4922
rect 6348 4870 6378 4922
rect 6402 4870 6412 4922
rect 6412 4870 6458 4922
rect 6482 4870 6528 4922
rect 6528 4870 6538 4922
rect 6562 4870 6592 4922
rect 6592 4870 6618 4922
rect 6322 4868 6378 4870
rect 6402 4868 6458 4870
rect 6482 4868 6538 4870
rect 6562 4868 6618 4870
rect 5249 4378 5305 4380
rect 5329 4378 5385 4380
rect 5409 4378 5465 4380
rect 5489 4378 5545 4380
rect 5249 4326 5275 4378
rect 5275 4326 5305 4378
rect 5329 4326 5339 4378
rect 5339 4326 5385 4378
rect 5409 4326 5455 4378
rect 5455 4326 5465 4378
rect 5489 4326 5519 4378
rect 5519 4326 5545 4378
rect 5249 4324 5305 4326
rect 5329 4324 5385 4326
rect 5409 4324 5465 4326
rect 5489 4324 5545 4326
rect 6734 4428 6736 4448
rect 6736 4428 6788 4448
rect 6788 4428 6790 4448
rect 6734 4392 6790 4428
rect 6322 3834 6378 3836
rect 6402 3834 6458 3836
rect 6482 3834 6538 3836
rect 6562 3834 6618 3836
rect 6322 3782 6348 3834
rect 6348 3782 6378 3834
rect 6402 3782 6412 3834
rect 6412 3782 6458 3834
rect 6482 3782 6528 3834
rect 6528 3782 6538 3834
rect 6562 3782 6592 3834
rect 6592 3782 6618 3834
rect 6322 3780 6378 3782
rect 6402 3780 6458 3782
rect 6482 3780 6538 3782
rect 6562 3780 6618 3782
rect 5249 3290 5305 3292
rect 5329 3290 5385 3292
rect 5409 3290 5465 3292
rect 5489 3290 5545 3292
rect 5249 3238 5275 3290
rect 5275 3238 5305 3290
rect 5329 3238 5339 3290
rect 5339 3238 5385 3290
rect 5409 3238 5455 3290
rect 5455 3238 5465 3290
rect 5489 3238 5519 3290
rect 5519 3238 5545 3290
rect 5249 3236 5305 3238
rect 5329 3236 5385 3238
rect 5409 3236 5465 3238
rect 5489 3236 5545 3238
rect 6322 2746 6378 2748
rect 6402 2746 6458 2748
rect 6482 2746 6538 2748
rect 6562 2746 6618 2748
rect 6322 2694 6348 2746
rect 6348 2694 6378 2746
rect 6402 2694 6412 2746
rect 6412 2694 6458 2746
rect 6482 2694 6528 2746
rect 6528 2694 6538 2746
rect 6562 2694 6592 2746
rect 6592 2694 6618 2746
rect 6322 2692 6378 2694
rect 6402 2692 6458 2694
rect 6482 2692 6538 2694
rect 6562 2692 6618 2694
rect 3102 2202 3158 2204
rect 3182 2202 3238 2204
rect 3262 2202 3318 2204
rect 3342 2202 3398 2204
rect 3102 2150 3128 2202
rect 3128 2150 3158 2202
rect 3182 2150 3192 2202
rect 3192 2150 3238 2202
rect 3262 2150 3308 2202
rect 3308 2150 3318 2202
rect 3342 2150 3372 2202
rect 3372 2150 3398 2202
rect 3102 2148 3158 2150
rect 3182 2148 3238 2150
rect 3262 2148 3318 2150
rect 3342 2148 3398 2150
rect 5249 2202 5305 2204
rect 5329 2202 5385 2204
rect 5409 2202 5465 2204
rect 5489 2202 5545 2204
rect 5249 2150 5275 2202
rect 5275 2150 5305 2202
rect 5329 2150 5339 2202
rect 5339 2150 5385 2202
rect 5409 2150 5455 2202
rect 5455 2150 5465 2202
rect 5489 2150 5519 2202
rect 5519 2150 5545 2202
rect 5249 2148 5305 2150
rect 5329 2148 5385 2150
rect 5409 2148 5465 2150
rect 5489 2148 5545 2150
rect 6826 40 6882 96
<< metal3 >>
rect 6821 8802 6887 8805
rect 7930 8802 8730 8832
rect 6821 8800 8730 8802
rect 6821 8744 6826 8800
rect 6882 8744 8730 8800
rect 6821 8742 8730 8744
rect 6821 8739 6887 8742
rect 7930 8712 8730 8742
rect 0 8530 800 8560
rect 1393 8530 1459 8533
rect 0 8528 1459 8530
rect 0 8472 1398 8528
rect 1454 8472 1459 8528
rect 0 8470 1459 8472
rect 0 8440 800 8470
rect 1393 8467 1459 8470
rect 2017 8192 2337 8193
rect 2017 8128 2025 8192
rect 2089 8128 2105 8192
rect 2169 8128 2185 8192
rect 2249 8128 2265 8192
rect 2329 8128 2337 8192
rect 2017 8127 2337 8128
rect 4164 8192 4484 8193
rect 4164 8128 4172 8192
rect 4236 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4484 8192
rect 4164 8127 4484 8128
rect 6310 8192 6630 8193
rect 6310 8128 6318 8192
rect 6382 8128 6398 8192
rect 6462 8128 6478 8192
rect 6542 8128 6558 8192
rect 6622 8128 6630 8192
rect 6310 8127 6630 8128
rect 3090 7648 3410 7649
rect 3090 7584 3098 7648
rect 3162 7584 3178 7648
rect 3242 7584 3258 7648
rect 3322 7584 3338 7648
rect 3402 7584 3410 7648
rect 3090 7583 3410 7584
rect 5237 7648 5557 7649
rect 5237 7584 5245 7648
rect 5309 7584 5325 7648
rect 5389 7584 5405 7648
rect 5469 7584 5485 7648
rect 5549 7584 5557 7648
rect 5237 7583 5557 7584
rect 2017 7104 2337 7105
rect 2017 7040 2025 7104
rect 2089 7040 2105 7104
rect 2169 7040 2185 7104
rect 2249 7040 2265 7104
rect 2329 7040 2337 7104
rect 2017 7039 2337 7040
rect 4164 7104 4484 7105
rect 4164 7040 4172 7104
rect 4236 7040 4252 7104
rect 4316 7040 4332 7104
rect 4396 7040 4412 7104
rect 4476 7040 4484 7104
rect 4164 7039 4484 7040
rect 6310 7104 6630 7105
rect 6310 7040 6318 7104
rect 6382 7040 6398 7104
rect 6462 7040 6478 7104
rect 6542 7040 6558 7104
rect 6622 7040 6630 7104
rect 6310 7039 6630 7040
rect 3090 6560 3410 6561
rect 3090 6496 3098 6560
rect 3162 6496 3178 6560
rect 3242 6496 3258 6560
rect 3322 6496 3338 6560
rect 3402 6496 3410 6560
rect 3090 6495 3410 6496
rect 5237 6560 5557 6561
rect 5237 6496 5245 6560
rect 5309 6496 5325 6560
rect 5389 6496 5405 6560
rect 5469 6496 5485 6560
rect 5549 6496 5557 6560
rect 5237 6495 5557 6496
rect 2017 6016 2337 6017
rect 2017 5952 2025 6016
rect 2089 5952 2105 6016
rect 2169 5952 2185 6016
rect 2249 5952 2265 6016
rect 2329 5952 2337 6016
rect 2017 5951 2337 5952
rect 4164 6016 4484 6017
rect 4164 5952 4172 6016
rect 4236 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4484 6016
rect 4164 5951 4484 5952
rect 6310 6016 6630 6017
rect 6310 5952 6318 6016
rect 6382 5952 6398 6016
rect 6462 5952 6478 6016
rect 6542 5952 6558 6016
rect 6622 5952 6630 6016
rect 6310 5951 6630 5952
rect 3090 5472 3410 5473
rect 3090 5408 3098 5472
rect 3162 5408 3178 5472
rect 3242 5408 3258 5472
rect 3322 5408 3338 5472
rect 3402 5408 3410 5472
rect 3090 5407 3410 5408
rect 5237 5472 5557 5473
rect 5237 5408 5245 5472
rect 5309 5408 5325 5472
rect 5389 5408 5405 5472
rect 5469 5408 5485 5472
rect 5549 5408 5557 5472
rect 5237 5407 5557 5408
rect 2017 4928 2337 4929
rect 2017 4864 2025 4928
rect 2089 4864 2105 4928
rect 2169 4864 2185 4928
rect 2249 4864 2265 4928
rect 2329 4864 2337 4928
rect 2017 4863 2337 4864
rect 4164 4928 4484 4929
rect 4164 4864 4172 4928
rect 4236 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4484 4928
rect 4164 4863 4484 4864
rect 6310 4928 6630 4929
rect 6310 4864 6318 4928
rect 6382 4864 6398 4928
rect 6462 4864 6478 4928
rect 6542 4864 6558 4928
rect 6622 4864 6630 4928
rect 6310 4863 6630 4864
rect 6729 4450 6795 4453
rect 7930 4450 8730 4480
rect 6729 4448 8730 4450
rect 6729 4392 6734 4448
rect 6790 4392 8730 4448
rect 6729 4390 8730 4392
rect 6729 4387 6795 4390
rect 3090 4384 3410 4385
rect 3090 4320 3098 4384
rect 3162 4320 3178 4384
rect 3242 4320 3258 4384
rect 3322 4320 3338 4384
rect 3402 4320 3410 4384
rect 3090 4319 3410 4320
rect 5237 4384 5557 4385
rect 5237 4320 5245 4384
rect 5309 4320 5325 4384
rect 5389 4320 5405 4384
rect 5469 4320 5485 4384
rect 5549 4320 5557 4384
rect 7930 4360 8730 4390
rect 5237 4319 5557 4320
rect 0 4178 800 4208
rect 1393 4178 1459 4181
rect 0 4176 1459 4178
rect 0 4120 1398 4176
rect 1454 4120 1459 4176
rect 0 4118 1459 4120
rect 0 4088 800 4118
rect 1393 4115 1459 4118
rect 2017 3840 2337 3841
rect 2017 3776 2025 3840
rect 2089 3776 2105 3840
rect 2169 3776 2185 3840
rect 2249 3776 2265 3840
rect 2329 3776 2337 3840
rect 2017 3775 2337 3776
rect 4164 3840 4484 3841
rect 4164 3776 4172 3840
rect 4236 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4484 3840
rect 4164 3775 4484 3776
rect 6310 3840 6630 3841
rect 6310 3776 6318 3840
rect 6382 3776 6398 3840
rect 6462 3776 6478 3840
rect 6542 3776 6558 3840
rect 6622 3776 6630 3840
rect 6310 3775 6630 3776
rect 3090 3296 3410 3297
rect 3090 3232 3098 3296
rect 3162 3232 3178 3296
rect 3242 3232 3258 3296
rect 3322 3232 3338 3296
rect 3402 3232 3410 3296
rect 3090 3231 3410 3232
rect 5237 3296 5557 3297
rect 5237 3232 5245 3296
rect 5309 3232 5325 3296
rect 5389 3232 5405 3296
rect 5469 3232 5485 3296
rect 5549 3232 5557 3296
rect 5237 3231 5557 3232
rect 2017 2752 2337 2753
rect 2017 2688 2025 2752
rect 2089 2688 2105 2752
rect 2169 2688 2185 2752
rect 2249 2688 2265 2752
rect 2329 2688 2337 2752
rect 2017 2687 2337 2688
rect 4164 2752 4484 2753
rect 4164 2688 4172 2752
rect 4236 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4484 2752
rect 4164 2687 4484 2688
rect 6310 2752 6630 2753
rect 6310 2688 6318 2752
rect 6382 2688 6398 2752
rect 6462 2688 6478 2752
rect 6542 2688 6558 2752
rect 6622 2688 6630 2752
rect 6310 2687 6630 2688
rect 3090 2208 3410 2209
rect 3090 2144 3098 2208
rect 3162 2144 3178 2208
rect 3242 2144 3258 2208
rect 3322 2144 3338 2208
rect 3402 2144 3410 2208
rect 3090 2143 3410 2144
rect 5237 2208 5557 2209
rect 5237 2144 5245 2208
rect 5309 2144 5325 2208
rect 5389 2144 5405 2208
rect 5469 2144 5485 2208
rect 5549 2144 5557 2208
rect 5237 2143 5557 2144
rect 6821 98 6887 101
rect 7930 98 8730 128
rect 6821 96 8730 98
rect 6821 40 6826 96
rect 6882 40 8730 96
rect 6821 38 8730 40
rect 6821 35 6887 38
rect 7930 8 8730 38
<< via3 >>
rect 2025 8188 2089 8192
rect 2025 8132 2029 8188
rect 2029 8132 2085 8188
rect 2085 8132 2089 8188
rect 2025 8128 2089 8132
rect 2105 8188 2169 8192
rect 2105 8132 2109 8188
rect 2109 8132 2165 8188
rect 2165 8132 2169 8188
rect 2105 8128 2169 8132
rect 2185 8188 2249 8192
rect 2185 8132 2189 8188
rect 2189 8132 2245 8188
rect 2245 8132 2249 8188
rect 2185 8128 2249 8132
rect 2265 8188 2329 8192
rect 2265 8132 2269 8188
rect 2269 8132 2325 8188
rect 2325 8132 2329 8188
rect 2265 8128 2329 8132
rect 4172 8188 4236 8192
rect 4172 8132 4176 8188
rect 4176 8132 4232 8188
rect 4232 8132 4236 8188
rect 4172 8128 4236 8132
rect 4252 8188 4316 8192
rect 4252 8132 4256 8188
rect 4256 8132 4312 8188
rect 4312 8132 4316 8188
rect 4252 8128 4316 8132
rect 4332 8188 4396 8192
rect 4332 8132 4336 8188
rect 4336 8132 4392 8188
rect 4392 8132 4396 8188
rect 4332 8128 4396 8132
rect 4412 8188 4476 8192
rect 4412 8132 4416 8188
rect 4416 8132 4472 8188
rect 4472 8132 4476 8188
rect 4412 8128 4476 8132
rect 6318 8188 6382 8192
rect 6318 8132 6322 8188
rect 6322 8132 6378 8188
rect 6378 8132 6382 8188
rect 6318 8128 6382 8132
rect 6398 8188 6462 8192
rect 6398 8132 6402 8188
rect 6402 8132 6458 8188
rect 6458 8132 6462 8188
rect 6398 8128 6462 8132
rect 6478 8188 6542 8192
rect 6478 8132 6482 8188
rect 6482 8132 6538 8188
rect 6538 8132 6542 8188
rect 6478 8128 6542 8132
rect 6558 8188 6622 8192
rect 6558 8132 6562 8188
rect 6562 8132 6618 8188
rect 6618 8132 6622 8188
rect 6558 8128 6622 8132
rect 3098 7644 3162 7648
rect 3098 7588 3102 7644
rect 3102 7588 3158 7644
rect 3158 7588 3162 7644
rect 3098 7584 3162 7588
rect 3178 7644 3242 7648
rect 3178 7588 3182 7644
rect 3182 7588 3238 7644
rect 3238 7588 3242 7644
rect 3178 7584 3242 7588
rect 3258 7644 3322 7648
rect 3258 7588 3262 7644
rect 3262 7588 3318 7644
rect 3318 7588 3322 7644
rect 3258 7584 3322 7588
rect 3338 7644 3402 7648
rect 3338 7588 3342 7644
rect 3342 7588 3398 7644
rect 3398 7588 3402 7644
rect 3338 7584 3402 7588
rect 5245 7644 5309 7648
rect 5245 7588 5249 7644
rect 5249 7588 5305 7644
rect 5305 7588 5309 7644
rect 5245 7584 5309 7588
rect 5325 7644 5389 7648
rect 5325 7588 5329 7644
rect 5329 7588 5385 7644
rect 5385 7588 5389 7644
rect 5325 7584 5389 7588
rect 5405 7644 5469 7648
rect 5405 7588 5409 7644
rect 5409 7588 5465 7644
rect 5465 7588 5469 7644
rect 5405 7584 5469 7588
rect 5485 7644 5549 7648
rect 5485 7588 5489 7644
rect 5489 7588 5545 7644
rect 5545 7588 5549 7644
rect 5485 7584 5549 7588
rect 2025 7100 2089 7104
rect 2025 7044 2029 7100
rect 2029 7044 2085 7100
rect 2085 7044 2089 7100
rect 2025 7040 2089 7044
rect 2105 7100 2169 7104
rect 2105 7044 2109 7100
rect 2109 7044 2165 7100
rect 2165 7044 2169 7100
rect 2105 7040 2169 7044
rect 2185 7100 2249 7104
rect 2185 7044 2189 7100
rect 2189 7044 2245 7100
rect 2245 7044 2249 7100
rect 2185 7040 2249 7044
rect 2265 7100 2329 7104
rect 2265 7044 2269 7100
rect 2269 7044 2325 7100
rect 2325 7044 2329 7100
rect 2265 7040 2329 7044
rect 4172 7100 4236 7104
rect 4172 7044 4176 7100
rect 4176 7044 4232 7100
rect 4232 7044 4236 7100
rect 4172 7040 4236 7044
rect 4252 7100 4316 7104
rect 4252 7044 4256 7100
rect 4256 7044 4312 7100
rect 4312 7044 4316 7100
rect 4252 7040 4316 7044
rect 4332 7100 4396 7104
rect 4332 7044 4336 7100
rect 4336 7044 4392 7100
rect 4392 7044 4396 7100
rect 4332 7040 4396 7044
rect 4412 7100 4476 7104
rect 4412 7044 4416 7100
rect 4416 7044 4472 7100
rect 4472 7044 4476 7100
rect 4412 7040 4476 7044
rect 6318 7100 6382 7104
rect 6318 7044 6322 7100
rect 6322 7044 6378 7100
rect 6378 7044 6382 7100
rect 6318 7040 6382 7044
rect 6398 7100 6462 7104
rect 6398 7044 6402 7100
rect 6402 7044 6458 7100
rect 6458 7044 6462 7100
rect 6398 7040 6462 7044
rect 6478 7100 6542 7104
rect 6478 7044 6482 7100
rect 6482 7044 6538 7100
rect 6538 7044 6542 7100
rect 6478 7040 6542 7044
rect 6558 7100 6622 7104
rect 6558 7044 6562 7100
rect 6562 7044 6618 7100
rect 6618 7044 6622 7100
rect 6558 7040 6622 7044
rect 3098 6556 3162 6560
rect 3098 6500 3102 6556
rect 3102 6500 3158 6556
rect 3158 6500 3162 6556
rect 3098 6496 3162 6500
rect 3178 6556 3242 6560
rect 3178 6500 3182 6556
rect 3182 6500 3238 6556
rect 3238 6500 3242 6556
rect 3178 6496 3242 6500
rect 3258 6556 3322 6560
rect 3258 6500 3262 6556
rect 3262 6500 3318 6556
rect 3318 6500 3322 6556
rect 3258 6496 3322 6500
rect 3338 6556 3402 6560
rect 3338 6500 3342 6556
rect 3342 6500 3398 6556
rect 3398 6500 3402 6556
rect 3338 6496 3402 6500
rect 5245 6556 5309 6560
rect 5245 6500 5249 6556
rect 5249 6500 5305 6556
rect 5305 6500 5309 6556
rect 5245 6496 5309 6500
rect 5325 6556 5389 6560
rect 5325 6500 5329 6556
rect 5329 6500 5385 6556
rect 5385 6500 5389 6556
rect 5325 6496 5389 6500
rect 5405 6556 5469 6560
rect 5405 6500 5409 6556
rect 5409 6500 5465 6556
rect 5465 6500 5469 6556
rect 5405 6496 5469 6500
rect 5485 6556 5549 6560
rect 5485 6500 5489 6556
rect 5489 6500 5545 6556
rect 5545 6500 5549 6556
rect 5485 6496 5549 6500
rect 2025 6012 2089 6016
rect 2025 5956 2029 6012
rect 2029 5956 2085 6012
rect 2085 5956 2089 6012
rect 2025 5952 2089 5956
rect 2105 6012 2169 6016
rect 2105 5956 2109 6012
rect 2109 5956 2165 6012
rect 2165 5956 2169 6012
rect 2105 5952 2169 5956
rect 2185 6012 2249 6016
rect 2185 5956 2189 6012
rect 2189 5956 2245 6012
rect 2245 5956 2249 6012
rect 2185 5952 2249 5956
rect 2265 6012 2329 6016
rect 2265 5956 2269 6012
rect 2269 5956 2325 6012
rect 2325 5956 2329 6012
rect 2265 5952 2329 5956
rect 4172 6012 4236 6016
rect 4172 5956 4176 6012
rect 4176 5956 4232 6012
rect 4232 5956 4236 6012
rect 4172 5952 4236 5956
rect 4252 6012 4316 6016
rect 4252 5956 4256 6012
rect 4256 5956 4312 6012
rect 4312 5956 4316 6012
rect 4252 5952 4316 5956
rect 4332 6012 4396 6016
rect 4332 5956 4336 6012
rect 4336 5956 4392 6012
rect 4392 5956 4396 6012
rect 4332 5952 4396 5956
rect 4412 6012 4476 6016
rect 4412 5956 4416 6012
rect 4416 5956 4472 6012
rect 4472 5956 4476 6012
rect 4412 5952 4476 5956
rect 6318 6012 6382 6016
rect 6318 5956 6322 6012
rect 6322 5956 6378 6012
rect 6378 5956 6382 6012
rect 6318 5952 6382 5956
rect 6398 6012 6462 6016
rect 6398 5956 6402 6012
rect 6402 5956 6458 6012
rect 6458 5956 6462 6012
rect 6398 5952 6462 5956
rect 6478 6012 6542 6016
rect 6478 5956 6482 6012
rect 6482 5956 6538 6012
rect 6538 5956 6542 6012
rect 6478 5952 6542 5956
rect 6558 6012 6622 6016
rect 6558 5956 6562 6012
rect 6562 5956 6618 6012
rect 6618 5956 6622 6012
rect 6558 5952 6622 5956
rect 3098 5468 3162 5472
rect 3098 5412 3102 5468
rect 3102 5412 3158 5468
rect 3158 5412 3162 5468
rect 3098 5408 3162 5412
rect 3178 5468 3242 5472
rect 3178 5412 3182 5468
rect 3182 5412 3238 5468
rect 3238 5412 3242 5468
rect 3178 5408 3242 5412
rect 3258 5468 3322 5472
rect 3258 5412 3262 5468
rect 3262 5412 3318 5468
rect 3318 5412 3322 5468
rect 3258 5408 3322 5412
rect 3338 5468 3402 5472
rect 3338 5412 3342 5468
rect 3342 5412 3398 5468
rect 3398 5412 3402 5468
rect 3338 5408 3402 5412
rect 5245 5468 5309 5472
rect 5245 5412 5249 5468
rect 5249 5412 5305 5468
rect 5305 5412 5309 5468
rect 5245 5408 5309 5412
rect 5325 5468 5389 5472
rect 5325 5412 5329 5468
rect 5329 5412 5385 5468
rect 5385 5412 5389 5468
rect 5325 5408 5389 5412
rect 5405 5468 5469 5472
rect 5405 5412 5409 5468
rect 5409 5412 5465 5468
rect 5465 5412 5469 5468
rect 5405 5408 5469 5412
rect 5485 5468 5549 5472
rect 5485 5412 5489 5468
rect 5489 5412 5545 5468
rect 5545 5412 5549 5468
rect 5485 5408 5549 5412
rect 2025 4924 2089 4928
rect 2025 4868 2029 4924
rect 2029 4868 2085 4924
rect 2085 4868 2089 4924
rect 2025 4864 2089 4868
rect 2105 4924 2169 4928
rect 2105 4868 2109 4924
rect 2109 4868 2165 4924
rect 2165 4868 2169 4924
rect 2105 4864 2169 4868
rect 2185 4924 2249 4928
rect 2185 4868 2189 4924
rect 2189 4868 2245 4924
rect 2245 4868 2249 4924
rect 2185 4864 2249 4868
rect 2265 4924 2329 4928
rect 2265 4868 2269 4924
rect 2269 4868 2325 4924
rect 2325 4868 2329 4924
rect 2265 4864 2329 4868
rect 4172 4924 4236 4928
rect 4172 4868 4176 4924
rect 4176 4868 4232 4924
rect 4232 4868 4236 4924
rect 4172 4864 4236 4868
rect 4252 4924 4316 4928
rect 4252 4868 4256 4924
rect 4256 4868 4312 4924
rect 4312 4868 4316 4924
rect 4252 4864 4316 4868
rect 4332 4924 4396 4928
rect 4332 4868 4336 4924
rect 4336 4868 4392 4924
rect 4392 4868 4396 4924
rect 4332 4864 4396 4868
rect 4412 4924 4476 4928
rect 4412 4868 4416 4924
rect 4416 4868 4472 4924
rect 4472 4868 4476 4924
rect 4412 4864 4476 4868
rect 6318 4924 6382 4928
rect 6318 4868 6322 4924
rect 6322 4868 6378 4924
rect 6378 4868 6382 4924
rect 6318 4864 6382 4868
rect 6398 4924 6462 4928
rect 6398 4868 6402 4924
rect 6402 4868 6458 4924
rect 6458 4868 6462 4924
rect 6398 4864 6462 4868
rect 6478 4924 6542 4928
rect 6478 4868 6482 4924
rect 6482 4868 6538 4924
rect 6538 4868 6542 4924
rect 6478 4864 6542 4868
rect 6558 4924 6622 4928
rect 6558 4868 6562 4924
rect 6562 4868 6618 4924
rect 6618 4868 6622 4924
rect 6558 4864 6622 4868
rect 3098 4380 3162 4384
rect 3098 4324 3102 4380
rect 3102 4324 3158 4380
rect 3158 4324 3162 4380
rect 3098 4320 3162 4324
rect 3178 4380 3242 4384
rect 3178 4324 3182 4380
rect 3182 4324 3238 4380
rect 3238 4324 3242 4380
rect 3178 4320 3242 4324
rect 3258 4380 3322 4384
rect 3258 4324 3262 4380
rect 3262 4324 3318 4380
rect 3318 4324 3322 4380
rect 3258 4320 3322 4324
rect 3338 4380 3402 4384
rect 3338 4324 3342 4380
rect 3342 4324 3398 4380
rect 3398 4324 3402 4380
rect 3338 4320 3402 4324
rect 5245 4380 5309 4384
rect 5245 4324 5249 4380
rect 5249 4324 5305 4380
rect 5305 4324 5309 4380
rect 5245 4320 5309 4324
rect 5325 4380 5389 4384
rect 5325 4324 5329 4380
rect 5329 4324 5385 4380
rect 5385 4324 5389 4380
rect 5325 4320 5389 4324
rect 5405 4380 5469 4384
rect 5405 4324 5409 4380
rect 5409 4324 5465 4380
rect 5465 4324 5469 4380
rect 5405 4320 5469 4324
rect 5485 4380 5549 4384
rect 5485 4324 5489 4380
rect 5489 4324 5545 4380
rect 5545 4324 5549 4380
rect 5485 4320 5549 4324
rect 2025 3836 2089 3840
rect 2025 3780 2029 3836
rect 2029 3780 2085 3836
rect 2085 3780 2089 3836
rect 2025 3776 2089 3780
rect 2105 3836 2169 3840
rect 2105 3780 2109 3836
rect 2109 3780 2165 3836
rect 2165 3780 2169 3836
rect 2105 3776 2169 3780
rect 2185 3836 2249 3840
rect 2185 3780 2189 3836
rect 2189 3780 2245 3836
rect 2245 3780 2249 3836
rect 2185 3776 2249 3780
rect 2265 3836 2329 3840
rect 2265 3780 2269 3836
rect 2269 3780 2325 3836
rect 2325 3780 2329 3836
rect 2265 3776 2329 3780
rect 4172 3836 4236 3840
rect 4172 3780 4176 3836
rect 4176 3780 4232 3836
rect 4232 3780 4236 3836
rect 4172 3776 4236 3780
rect 4252 3836 4316 3840
rect 4252 3780 4256 3836
rect 4256 3780 4312 3836
rect 4312 3780 4316 3836
rect 4252 3776 4316 3780
rect 4332 3836 4396 3840
rect 4332 3780 4336 3836
rect 4336 3780 4392 3836
rect 4392 3780 4396 3836
rect 4332 3776 4396 3780
rect 4412 3836 4476 3840
rect 4412 3780 4416 3836
rect 4416 3780 4472 3836
rect 4472 3780 4476 3836
rect 4412 3776 4476 3780
rect 6318 3836 6382 3840
rect 6318 3780 6322 3836
rect 6322 3780 6378 3836
rect 6378 3780 6382 3836
rect 6318 3776 6382 3780
rect 6398 3836 6462 3840
rect 6398 3780 6402 3836
rect 6402 3780 6458 3836
rect 6458 3780 6462 3836
rect 6398 3776 6462 3780
rect 6478 3836 6542 3840
rect 6478 3780 6482 3836
rect 6482 3780 6538 3836
rect 6538 3780 6542 3836
rect 6478 3776 6542 3780
rect 6558 3836 6622 3840
rect 6558 3780 6562 3836
rect 6562 3780 6618 3836
rect 6618 3780 6622 3836
rect 6558 3776 6622 3780
rect 3098 3292 3162 3296
rect 3098 3236 3102 3292
rect 3102 3236 3158 3292
rect 3158 3236 3162 3292
rect 3098 3232 3162 3236
rect 3178 3292 3242 3296
rect 3178 3236 3182 3292
rect 3182 3236 3238 3292
rect 3238 3236 3242 3292
rect 3178 3232 3242 3236
rect 3258 3292 3322 3296
rect 3258 3236 3262 3292
rect 3262 3236 3318 3292
rect 3318 3236 3322 3292
rect 3258 3232 3322 3236
rect 3338 3292 3402 3296
rect 3338 3236 3342 3292
rect 3342 3236 3398 3292
rect 3398 3236 3402 3292
rect 3338 3232 3402 3236
rect 5245 3292 5309 3296
rect 5245 3236 5249 3292
rect 5249 3236 5305 3292
rect 5305 3236 5309 3292
rect 5245 3232 5309 3236
rect 5325 3292 5389 3296
rect 5325 3236 5329 3292
rect 5329 3236 5385 3292
rect 5385 3236 5389 3292
rect 5325 3232 5389 3236
rect 5405 3292 5469 3296
rect 5405 3236 5409 3292
rect 5409 3236 5465 3292
rect 5465 3236 5469 3292
rect 5405 3232 5469 3236
rect 5485 3292 5549 3296
rect 5485 3236 5489 3292
rect 5489 3236 5545 3292
rect 5545 3236 5549 3292
rect 5485 3232 5549 3236
rect 2025 2748 2089 2752
rect 2025 2692 2029 2748
rect 2029 2692 2085 2748
rect 2085 2692 2089 2748
rect 2025 2688 2089 2692
rect 2105 2748 2169 2752
rect 2105 2692 2109 2748
rect 2109 2692 2165 2748
rect 2165 2692 2169 2748
rect 2105 2688 2169 2692
rect 2185 2748 2249 2752
rect 2185 2692 2189 2748
rect 2189 2692 2245 2748
rect 2245 2692 2249 2748
rect 2185 2688 2249 2692
rect 2265 2748 2329 2752
rect 2265 2692 2269 2748
rect 2269 2692 2325 2748
rect 2325 2692 2329 2748
rect 2265 2688 2329 2692
rect 4172 2748 4236 2752
rect 4172 2692 4176 2748
rect 4176 2692 4232 2748
rect 4232 2692 4236 2748
rect 4172 2688 4236 2692
rect 4252 2748 4316 2752
rect 4252 2692 4256 2748
rect 4256 2692 4312 2748
rect 4312 2692 4316 2748
rect 4252 2688 4316 2692
rect 4332 2748 4396 2752
rect 4332 2692 4336 2748
rect 4336 2692 4392 2748
rect 4392 2692 4396 2748
rect 4332 2688 4396 2692
rect 4412 2748 4476 2752
rect 4412 2692 4416 2748
rect 4416 2692 4472 2748
rect 4472 2692 4476 2748
rect 4412 2688 4476 2692
rect 6318 2748 6382 2752
rect 6318 2692 6322 2748
rect 6322 2692 6378 2748
rect 6378 2692 6382 2748
rect 6318 2688 6382 2692
rect 6398 2748 6462 2752
rect 6398 2692 6402 2748
rect 6402 2692 6458 2748
rect 6458 2692 6462 2748
rect 6398 2688 6462 2692
rect 6478 2748 6542 2752
rect 6478 2692 6482 2748
rect 6482 2692 6538 2748
rect 6538 2692 6542 2748
rect 6478 2688 6542 2692
rect 6558 2748 6622 2752
rect 6558 2692 6562 2748
rect 6562 2692 6618 2748
rect 6618 2692 6622 2748
rect 6558 2688 6622 2692
rect 3098 2204 3162 2208
rect 3098 2148 3102 2204
rect 3102 2148 3158 2204
rect 3158 2148 3162 2204
rect 3098 2144 3162 2148
rect 3178 2204 3242 2208
rect 3178 2148 3182 2204
rect 3182 2148 3238 2204
rect 3238 2148 3242 2204
rect 3178 2144 3242 2148
rect 3258 2204 3322 2208
rect 3258 2148 3262 2204
rect 3262 2148 3318 2204
rect 3318 2148 3322 2204
rect 3258 2144 3322 2148
rect 3338 2204 3402 2208
rect 3338 2148 3342 2204
rect 3342 2148 3398 2204
rect 3398 2148 3402 2204
rect 3338 2144 3402 2148
rect 5245 2204 5309 2208
rect 5245 2148 5249 2204
rect 5249 2148 5305 2204
rect 5305 2148 5309 2204
rect 5245 2144 5309 2148
rect 5325 2204 5389 2208
rect 5325 2148 5329 2204
rect 5329 2148 5385 2204
rect 5385 2148 5389 2204
rect 5325 2144 5389 2148
rect 5405 2204 5469 2208
rect 5405 2148 5409 2204
rect 5409 2148 5465 2204
rect 5465 2148 5469 2204
rect 5405 2144 5469 2148
rect 5485 2204 5549 2208
rect 5485 2148 5489 2204
rect 5489 2148 5545 2204
rect 5545 2148 5549 2204
rect 5485 2144 5549 2148
<< metal4 >>
rect 2017 8192 2337 8208
rect 2017 8128 2025 8192
rect 2089 8128 2105 8192
rect 2169 8128 2185 8192
rect 2249 8128 2265 8192
rect 2329 8128 2337 8192
rect 2017 7232 2337 8128
rect 2017 7104 2059 7232
rect 2295 7104 2337 7232
rect 2017 7040 2025 7104
rect 2329 7040 2337 7104
rect 2017 6996 2059 7040
rect 2295 6996 2337 7040
rect 2017 6016 2337 6996
rect 2017 5952 2025 6016
rect 2089 5952 2105 6016
rect 2169 5952 2185 6016
rect 2249 5952 2265 6016
rect 2329 5952 2337 6016
rect 2017 5238 2337 5952
rect 2017 5002 2059 5238
rect 2295 5002 2337 5238
rect 2017 4928 2337 5002
rect 2017 4864 2025 4928
rect 2089 4864 2105 4928
rect 2169 4864 2185 4928
rect 2249 4864 2265 4928
rect 2329 4864 2337 4928
rect 2017 3840 2337 4864
rect 2017 3776 2025 3840
rect 2089 3776 2105 3840
rect 2169 3776 2185 3840
rect 2249 3776 2265 3840
rect 2329 3776 2337 3840
rect 2017 3243 2337 3776
rect 2017 3007 2059 3243
rect 2295 3007 2337 3243
rect 2017 2752 2337 3007
rect 2017 2688 2025 2752
rect 2089 2688 2105 2752
rect 2169 2688 2185 2752
rect 2249 2688 2265 2752
rect 2329 2688 2337 2752
rect 2017 2128 2337 2688
rect 3090 7648 3410 8208
rect 3090 7584 3098 7648
rect 3162 7584 3178 7648
rect 3242 7584 3258 7648
rect 3322 7584 3338 7648
rect 3402 7584 3410 7648
rect 3090 6560 3410 7584
rect 3090 6496 3098 6560
rect 3162 6496 3178 6560
rect 3242 6496 3258 6560
rect 3322 6496 3338 6560
rect 3402 6496 3410 6560
rect 3090 6235 3410 6496
rect 3090 5999 3132 6235
rect 3368 5999 3410 6235
rect 3090 5472 3410 5999
rect 3090 5408 3098 5472
rect 3162 5408 3178 5472
rect 3242 5408 3258 5472
rect 3322 5408 3338 5472
rect 3402 5408 3410 5472
rect 3090 4384 3410 5408
rect 3090 4320 3098 4384
rect 3162 4320 3178 4384
rect 3242 4320 3258 4384
rect 3322 4320 3338 4384
rect 3402 4320 3410 4384
rect 3090 4240 3410 4320
rect 3090 4004 3132 4240
rect 3368 4004 3410 4240
rect 3090 3296 3410 4004
rect 3090 3232 3098 3296
rect 3162 3232 3178 3296
rect 3242 3232 3258 3296
rect 3322 3232 3338 3296
rect 3402 3232 3410 3296
rect 3090 2208 3410 3232
rect 3090 2144 3098 2208
rect 3162 2144 3178 2208
rect 3242 2144 3258 2208
rect 3322 2144 3338 2208
rect 3402 2144 3410 2208
rect 3090 2128 3410 2144
rect 4164 8192 4484 8208
rect 4164 8128 4172 8192
rect 4236 8128 4252 8192
rect 4316 8128 4332 8192
rect 4396 8128 4412 8192
rect 4476 8128 4484 8192
rect 4164 7232 4484 8128
rect 4164 7104 4206 7232
rect 4442 7104 4484 7232
rect 4164 7040 4172 7104
rect 4476 7040 4484 7104
rect 4164 6996 4206 7040
rect 4442 6996 4484 7040
rect 4164 6016 4484 6996
rect 4164 5952 4172 6016
rect 4236 5952 4252 6016
rect 4316 5952 4332 6016
rect 4396 5952 4412 6016
rect 4476 5952 4484 6016
rect 4164 5238 4484 5952
rect 4164 5002 4206 5238
rect 4442 5002 4484 5238
rect 4164 4928 4484 5002
rect 4164 4864 4172 4928
rect 4236 4864 4252 4928
rect 4316 4864 4332 4928
rect 4396 4864 4412 4928
rect 4476 4864 4484 4928
rect 4164 3840 4484 4864
rect 4164 3776 4172 3840
rect 4236 3776 4252 3840
rect 4316 3776 4332 3840
rect 4396 3776 4412 3840
rect 4476 3776 4484 3840
rect 4164 3243 4484 3776
rect 4164 3007 4206 3243
rect 4442 3007 4484 3243
rect 4164 2752 4484 3007
rect 4164 2688 4172 2752
rect 4236 2688 4252 2752
rect 4316 2688 4332 2752
rect 4396 2688 4412 2752
rect 4476 2688 4484 2752
rect 4164 2128 4484 2688
rect 5237 7648 5557 8208
rect 5237 7584 5245 7648
rect 5309 7584 5325 7648
rect 5389 7584 5405 7648
rect 5469 7584 5485 7648
rect 5549 7584 5557 7648
rect 5237 6560 5557 7584
rect 5237 6496 5245 6560
rect 5309 6496 5325 6560
rect 5389 6496 5405 6560
rect 5469 6496 5485 6560
rect 5549 6496 5557 6560
rect 5237 6235 5557 6496
rect 5237 5999 5279 6235
rect 5515 5999 5557 6235
rect 5237 5472 5557 5999
rect 5237 5408 5245 5472
rect 5309 5408 5325 5472
rect 5389 5408 5405 5472
rect 5469 5408 5485 5472
rect 5549 5408 5557 5472
rect 5237 4384 5557 5408
rect 5237 4320 5245 4384
rect 5309 4320 5325 4384
rect 5389 4320 5405 4384
rect 5469 4320 5485 4384
rect 5549 4320 5557 4384
rect 5237 4240 5557 4320
rect 5237 4004 5279 4240
rect 5515 4004 5557 4240
rect 5237 3296 5557 4004
rect 5237 3232 5245 3296
rect 5309 3232 5325 3296
rect 5389 3232 5405 3296
rect 5469 3232 5485 3296
rect 5549 3232 5557 3296
rect 5237 2208 5557 3232
rect 5237 2144 5245 2208
rect 5309 2144 5325 2208
rect 5389 2144 5405 2208
rect 5469 2144 5485 2208
rect 5549 2144 5557 2208
rect 5237 2128 5557 2144
rect 6310 8192 6630 8208
rect 6310 8128 6318 8192
rect 6382 8128 6398 8192
rect 6462 8128 6478 8192
rect 6542 8128 6558 8192
rect 6622 8128 6630 8192
rect 6310 7232 6630 8128
rect 6310 7104 6352 7232
rect 6588 7104 6630 7232
rect 6310 7040 6318 7104
rect 6622 7040 6630 7104
rect 6310 6996 6352 7040
rect 6588 6996 6630 7040
rect 6310 6016 6630 6996
rect 6310 5952 6318 6016
rect 6382 5952 6398 6016
rect 6462 5952 6478 6016
rect 6542 5952 6558 6016
rect 6622 5952 6630 6016
rect 6310 5238 6630 5952
rect 6310 5002 6352 5238
rect 6588 5002 6630 5238
rect 6310 4928 6630 5002
rect 6310 4864 6318 4928
rect 6382 4864 6398 4928
rect 6462 4864 6478 4928
rect 6542 4864 6558 4928
rect 6622 4864 6630 4928
rect 6310 3840 6630 4864
rect 6310 3776 6318 3840
rect 6382 3776 6398 3840
rect 6462 3776 6478 3840
rect 6542 3776 6558 3840
rect 6622 3776 6630 3840
rect 6310 3243 6630 3776
rect 6310 3007 6352 3243
rect 6588 3007 6630 3243
rect 6310 2752 6630 3007
rect 6310 2688 6318 2752
rect 6382 2688 6398 2752
rect 6462 2688 6478 2752
rect 6542 2688 6558 2752
rect 6622 2688 6630 2752
rect 6310 2128 6630 2688
<< via4 >>
rect 2059 7104 2295 7232
rect 2059 7040 2089 7104
rect 2089 7040 2105 7104
rect 2105 7040 2169 7104
rect 2169 7040 2185 7104
rect 2185 7040 2249 7104
rect 2249 7040 2265 7104
rect 2265 7040 2295 7104
rect 2059 6996 2295 7040
rect 2059 5002 2295 5238
rect 2059 3007 2295 3243
rect 3132 5999 3368 6235
rect 3132 4004 3368 4240
rect 4206 7104 4442 7232
rect 4206 7040 4236 7104
rect 4236 7040 4252 7104
rect 4252 7040 4316 7104
rect 4316 7040 4332 7104
rect 4332 7040 4396 7104
rect 4396 7040 4412 7104
rect 4412 7040 4442 7104
rect 4206 6996 4442 7040
rect 4206 5002 4442 5238
rect 4206 3007 4442 3243
rect 5279 5999 5515 6235
rect 5279 4004 5515 4240
rect 6352 7104 6588 7232
rect 6352 7040 6382 7104
rect 6382 7040 6398 7104
rect 6398 7040 6462 7104
rect 6462 7040 6478 7104
rect 6478 7040 6542 7104
rect 6542 7040 6558 7104
rect 6558 7040 6588 7104
rect 6352 6996 6588 7040
rect 6352 5002 6588 5238
rect 6352 3007 6588 3243
<< metal5 >>
rect 1104 7232 7544 7274
rect 1104 6996 2059 7232
rect 2295 6996 4206 7232
rect 4442 6996 6352 7232
rect 6588 6996 7544 7232
rect 1104 6954 7544 6996
rect 1104 6235 7544 6277
rect 1104 5999 3132 6235
rect 3368 5999 5279 6235
rect 5515 5999 7544 6235
rect 1104 5957 7544 5999
rect 1104 5238 7544 5280
rect 1104 5002 2059 5238
rect 2295 5002 4206 5238
rect 4442 5002 6352 5238
rect 6588 5002 7544 5238
rect 1104 4960 7544 5002
rect 1104 4240 7544 4282
rect 1104 4004 3132 4240
rect 3368 4004 5279 4240
rect 5515 4004 7544 4240
rect 1104 3962 7544 4004
rect 1104 3243 7544 3286
rect 1104 3007 2059 3243
rect 2295 3007 4206 3243
rect 4442 3007 6352 3243
rect 6588 3007 7544 3243
rect 1104 2965 7544 3007
use sky130_fd_sc_hd__decap_12  FILLER_0_6
timestamp 1629539722
transform 1 0 1656 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1629539722
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1629539722
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1629539722
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1629539722
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp 1629539722
transform 1 0 2760 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1629539722
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1629539722
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1629539722
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_29
timestamp 1629539722
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1629539722
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_22
timestamp 1629539722
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41
timestamp 1629539722
transform 1 0 4876 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1629539722
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 1629539722
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1629539722
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1629539722
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57
timestamp 1629539722
transform 1 0 6348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1629539722
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1629539722
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_57
timestamp 1629539722
transform 1 0 6348 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_23
timestamp 1629539722
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_24
timestamp 1629539722
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1629539722
transform 1 0 6624 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 1629539722
transform 1 0 7084 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1629539722
transform -1 0 7544 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1629539722
transform -1 0 7544 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1629539722
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1629539722
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1629539722
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1629539722
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1629539722
transform 1 0 4048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_25
timestamp 1629539722
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _17_
timestamp 1629539722
transform 1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_40
timestamp 1629539722
transform 1 0 4784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_45
timestamp 1629539722
transform 1 0 5244 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _12_
timestamp 1629539722
transform -1 0 5888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _14_
timestamp 1629539722
transform -1 0 5244 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_52
timestamp 1629539722
transform 1 0 5888 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_64
timestamp 1629539722
transform 1 0 6992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1629539722
transform -1 0 7544 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1629539722
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1629539722
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_15
timestamp 1629539722
transform 1 0 2484 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _20_
timestamp 1629539722
transform 1 0 3036 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_3_30
timestamp 1629539722
transform 1 0 3864 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_38
timestamp 1629539722
transform 1 0 4600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_47
timestamp 1629539722
transform 1 0 5428 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _16_
timestamp 1629539722
transform 1 0 4692 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1629539722
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_57
timestamp 1629539722
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_26
timestamp 1629539722
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_65
timestamp 1629539722
transform 1 0 7084 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1629539722
transform -1 0 7544 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_6
timestamp 1629539722
transform 1 0 1656 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1629539722
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1629539722
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1629539722
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _19_
timestamp 1629539722
transform 1 0 2760 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_36
timestamp 1629539722
transform 1 0 4416 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_27
timestamp 1629539722
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_1  _23_
timestamp 1629539722
transform 1 0 3772 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_4_40
timestamp 1629539722
transform 1 0 4784 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_50
timestamp 1629539722
transform 1 0 5704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _15_
timestamp 1629539722
transform -1 0 5704 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_4_58
timestamp 1629539722
transform 1 0 6440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_63
timestamp 1629539722
transform 1 0 6900 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  output11
timestamp 1629539722
transform 1 0 6532 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1629539722
transform -1 0 7544 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1629539722
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1629539722
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_15
timestamp 1629539722
transform 1 0 2484 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_23
timestamp 1629539722
transform 1 0 3220 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_1  _22_
timestamp 1629539722
transform -1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_28
timestamp 1629539722
transform 1 0 3680 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1629539722
transform 1 0 4324 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _21_
timestamp 1629539722
transform 1 0 4048 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_47
timestamp 1629539722
transform 1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _25_
timestamp 1629539722
transform -1 0 5428 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1629539722
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_60
timestamp 1629539722
transform 1 0 6624 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28
timestamp 1629539722
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _24_
timestamp 1629539722
transform 1 0 6348 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_66
timestamp 1629539722
transform 1 0 7176 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1629539722
transform -1 0 7544 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1629539722
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1629539722
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1629539722
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1629539722
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1629539722
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1629539722
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1629539722
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_32
timestamp 1629539722
transform 1 0 4048 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1629539722
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1629539722
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _18_
timestamp 1629539722
transform -1 0 4048 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 1629539722
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_39
timestamp 1629539722
transform 1 0 4692 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_48
timestamp 1629539722
transform 1 0 5520 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1629539722
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1629539722
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _13_
timestamp 1629539722
transform -1 0 5520 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_6_60
timestamp 1629539722
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1629539722
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1629539722
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1629539722
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_66
timestamp 1629539722
transform 1 0 7176 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_65
timestamp 1629539722
transform 1 0 7084 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1629539722
transform -1 0 7544 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1629539722
transform -1 0 7544 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1629539722
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1629539722
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1629539722
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1629539722
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1629539722
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1629539722
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1629539722
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1629539722
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_65
timestamp 1629539722
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1629539722
transform -1 0 7544 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_6
timestamp 1629539722
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1629539722
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 1629539722
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_18
timestamp 1629539722
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_30
timestamp 1629539722
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_42
timestamp 1629539722
transform 1 0 4968 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_54
timestamp 1629539722
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 1629539722
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_63
timestamp 1629539722
transform 1 0 6900 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1629539722
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1629539722
transform -1 0 6900 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1629539722
transform -1 0 7544 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_11
timestamp 1629539722
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1629539722
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1629539722
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  output9
timestamp 1629539722
transform -1 0 2116 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_23
timestamp 1629539722
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1629539722
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_29
timestamp 1629539722
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1629539722
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  output10
timestamp 1629539722
transform -1 0 4692 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_39
timestamp 1629539722
transform 1 0 4692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_51
timestamp 1629539722
transform 1 0 5796 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_55
timestamp 1629539722
transform 1 0 6164 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_57
timestamp 1629539722
transform 1 0 6348 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_63
timestamp 1629539722
transform 1 0 6900 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1629539722
transform 1 0 6256 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1629539722
transform -1 0 6900 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1629539722
transform -1 0 7544 0 1 7616
box -38 -48 314 592
<< labels >>
rlabel metal3 s 0 8440 800 8560 4 A_in[0]
port 1 nsew
rlabel metal3 s 7930 8 8730 128 4 A_in[1]
port 2 nsew
rlabel metal2 s 18 0 74 800 4 A_in[2]
port 3 nsew
rlabel metal2 s 7194 10074 7250 10874 4 A_in[3]
port 4 nsew
rlabel metal2 s 5906 0 5962 800 4 B_in[0]
port 5 nsew
rlabel metal3 s 0 4088 800 4208 4 B_in[1]
port 6 nsew
rlabel metal3 s 7930 8712 8730 8832 4 B_in[2]
port 7 nsew
rlabel metal2 s 2962 0 3018 800 4 B_in[3]
port 8 nsew
rlabel metal5 s 1104 3962 7544 4282 4 VGND
port 9 nsew
rlabel metal5 s 1104 2966 7544 3286 4 VPWR
port 10 nsew
rlabel metal2 s 1306 10074 1362 10874 4 equal_to
port 11 nsew
rlabel metal2 s 4250 10074 4306 10874 4 greater_than
port 12 nsew
rlabel metal3 s 7930 4360 8730 4480 4 less_than
port 13 nsew
<< properties >>
string FIXED_BBOX 0 0 8730 10874
<< end >>
