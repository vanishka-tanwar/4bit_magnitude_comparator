* SPICE3 file created from dvsd_cmp.ext - technology: sky130A

.subckt dvsd_cmp A_in[0] A_in[1] A_in[2] A_in[3] B_in[0] B_in[1] B_in[2] B_in[3] VGND
+ VPWR equal_to greater_than less_than
C0 _13_/Y _24_/Y 0.08fF
C1 B_in[1] _14_/A 0.02fF
C2 _26_/A _26_/Y 0.05fF
C3 _20_/B2 _14_/A 0.03fF
C4 _22_/A VPWR 2.90fF
C5 _26_/B _21_/A 0.11fF
C6 _26_/Y _24_/A 0.31fF
C7 _15_/X _14_/B 0.13fF
C8 _21_/Y VPWR 1.07fF
C9 _18_/Y VPWR 0.34fF
C10 A_in[2] _20_/B2 0.02fF
C11 B_in[1] VPWR 0.02fF
C12 _18_/A B_in[2] 0.02fF
C13 VPWR _18_/A 1.59fF
C14 _12_/A VPWR 1.32fF
C15 _22_/A _15_/X 0.09fF
C16 greater_than _26_/B 0.10fF
C17 _20_/B2 VPWR 1.78fF
C18 _19_/Y _14_/A 1.18fF
C19 _26_/A _26_/B 0.55fF
C20 _22_/A _22_/B 1.14fF
C21 _21_/A _14_/A 0.03fF
C22 _22_/Y _19_/Y 0.18fF
C23 _21_/A _22_/Y 0.22fF
C24 less_than VPWR 0.03fF
C25 _21_/Y _15_/X 0.05fF
C26 VPWR _24_/Y 0.81fF
C27 _13_/A _26_/B 0.14fF
C28 _22_/A _14_/B 0.01fF
C29 _13_/Y _26_/A 0.07fF
C30 _26_/B _24_/A 0.63fF
C31 _22_/B _18_/Y 0.49fF
C32 _17_/A VPWR 0.95fF
C33 _13_/A _13_/Y 0.51fF
C34 A_in[1] _12_/A 0.02fF
C35 A_in[0] _24_/A 0.02fF
C36 _13_/Y _24_/A 0.69fF
C37 _22_/B _20_/B2 0.18fF
C38 VPWR _19_/Y 0.36fF
C39 _26_/A _14_/A 0.58fF
C40 _21_/A VPWR 0.60fF
C41 _12_/A _14_/B 0.06fF
C42 _26_/A _22_/Y 0.05fF
C43 _15_/X _24_/Y 0.03fF
C44 _26_/B _26_/Y 2.14fF
C45 _21_/Y _22_/A 0.06fF
C46 _13_/A _14_/A 1.05fF
C47 _22_/A _18_/Y 1.41fF
C48 _26_/A _14_/Y 0.18fF
C49 _16_/X _14_/A 0.09fF
C50 _24_/A _14_/A 0.17fF
C51 _16_/X _22_/Y 0.04fF
C52 _22_/A _18_/A 0.05fF
C53 _17_/A B_in[3] 0.02fF
C54 _17_/A _22_/B 0.05fF
C55 _13_/A _14_/Y 0.07fF
C56 _22_/A _20_/B2 0.05fF
C57 greater_than VPWR 0.48fF
C58 _14_/Y _24_/A 0.04fF
C59 _15_/X _21_/A 0.03fF
C60 _26_/A VPWR 0.76fF
C61 _22_/B _19_/Y 1.27fF
C62 _18_/Y _18_/A 0.05fF
C63 _22_/B _21_/A 0.72fF
C64 _22_/A _24_/Y 0.16fF
C65 _26_/B equal_to 0.04fF
C66 _20_/B2 _18_/Y 0.29fF
C67 _13_/A VPWR 1.46fF
C68 equal_to A_in[0] 0.56fF
C69 _16_/X VPWR 0.29fF
C70 VPWR _24_/A 5.67fF
C71 B_in[0] VPWR 0.03fF
C72 _26_/A _15_/X 0.33fF
C73 _22_/A _19_/Y 0.74fF
C74 _22_/A _21_/A 1.18fF
C75 _13_/Y _26_/B 0.13fF
C76 _22_/B _26_/A 0.17fF
C77 _13_/A _15_/X 1.17fF
C78 _26_/Y VPWR 0.51fF
C79 _21_/Y _19_/Y 0.01fF
C80 _21_/Y _21_/A 0.24fF
C81 _16_/X _15_/X 0.02fF
C82 _26_/A _14_/B 0.27fF
C83 _18_/Y _19_/Y 0.69fF
C84 _15_/X _24_/A 0.73fF
C85 _18_/Y _21_/A 0.17fF
C86 _17_/A _20_/B2 0.01fF
C87 _16_/X _22_/B 0.01fF
C88 _13_/A _14_/B 0.35fF
C89 _16_/X _14_/B 0.00fF
C90 _20_/B2 _19_/Y 0.48fF
C91 _20_/B2 _21_/A 0.01fF
C92 _14_/B _24_/A 0.08fF
C93 _22_/A _26_/A 0.05fF
C94 A_in[3] B_in[2] 0.29fF
C95 _13_/Y _14_/A 0.01fF
C96 A_in[3] VPWR 0.17fF
C97 _13_/A _22_/A 0.16fF
C98 _21_/A _24_/Y 0.01fF
C99 equal_to VPWR 0.33fF
C100 _21_/Y _26_/A 0.29fF
C101 _13_/Y _14_/Y 0.01fF
C102 _26_/A _18_/Y 0.01fF
C103 _22_/A _24_/A 0.40fF
C104 _17_/A _21_/A 0.01fF
C105 _26_/B VPWR 1.06fF
C106 _26_/A _18_/A 0.15fF
C107 _16_/X _21_/Y 0.08fF
C108 _22_/Y _14_/A 0.18fF
C109 VPWR A_in[0] 0.11fF
C110 _21_/Y _24_/A 0.06fF
C111 _13_/A _18_/A 0.64fF
C112 _13_/Y VPWR 0.28fF
C113 _13_/A _12_/A 0.02fF
C114 _21_/A _19_/Y 0.05fF
C115 _14_/Y _14_/A 0.36fF
C116 less_than _26_/A 0.05fF
C117 _24_/A _18_/A 0.03fF
C118 _12_/A B_in[0] 0.04fF
C119 _26_/B _15_/X 0.05fF
C120 _13_/A _24_/Y 0.15fF
C121 VPWR _14_/A 1.72fF
C122 _24_/A _24_/Y 1.21fF
C123 VPWR _22_/Y 1.03fF
C124 _26_/Y _18_/A 0.16fF
C125 _13_/Y _15_/X 0.13fF
C126 _22_/A A_in[3] 0.02fF
C127 _26_/A _19_/Y 0.14fF
C128 _26_/A _21_/A 0.32fF
C129 _14_/Y VPWR 0.88fF
C130 A_in[2] VPWR 0.07fF
C131 _13_/A _21_/A 0.02fF
C132 _13_/Y _14_/B 0.36fF
C133 _16_/X _19_/Y 0.01fF
C134 _22_/A _26_/B 0.20fF
C135 _15_/X _14_/A 0.30fF
C136 VPWR B_in[2] 0.13fF
C137 _22_/B _14_/A 0.36fF
C138 _22_/B _22_/Y 0.37fF
C139 _22_/A _13_/Y 0.07fF
C140 _21_/Y _26_/B 0.02fF
C141 _14_/B _14_/A 1.35fF
C142 _26_/B _18_/A 0.36fF
C143 _13_/A _26_/A 0.23fF
C144 _16_/X _26_/A 0.24fF
C145 _14_/Y _14_/B 0.23fF
C146 _26_/A _24_/A 0.55fF
C147 _22_/A _14_/A 0.41fF
C148 _15_/X VPWR 0.38fF
C149 A_in[1] VPWR 0.02fF
C150 _13_/Y _18_/A 0.12fF
C151 B_in[3] VPWR 0.03fF
C152 _22_/A _22_/Y 0.36fF
C153 _22_/B VPWR 0.76fF
C154 _13_/A _24_/A 0.38fF
C155 _26_/B _24_/Y 0.45fF
C156 _21_/Y _14_/A 0.52fF
C157 _22_/A _14_/Y 0.02fF
C158 VPWR _14_/B 0.26fF
C159 _21_/Y _22_/Y 0.12fF
C160 _18_/Y _14_/A 0.14fF
C161 greater_than _26_/Y 0.08fF
C162 _13_/A B_in[0] 0.02fF
XFILLER_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput10 _26_/Y VGND VGND VPWR VPWR greater_than sky130_fd_sc_hd__clkbuf_2
XFILLER_3_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xoutput9 _26_/B VGND VGND VPWR VPWR equal_to sky130_fd_sc_hd__clkbuf_2
Xoutput11 _26_/A VGND VGND VPWR VPWR less_than sky130_fd_sc_hd__clkbuf_2
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_26_ _26_/A _26_/B VGND VGND VPWR VPWR _26_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_25_ _24_/Y _13_/A _15_/X _21_/A VGND VGND VPWR VPWR _26_/B sky130_fd_sc_hd__o211a_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_24_ _24_/A VGND VGND VPWR VPWR _24_/Y sky130_fd_sc_hd__inv_2
XFILLER_10_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_23_ _16_/X _21_/Y _19_/Y _22_/Y VGND VGND VPWR VPWR _26_/A sky130_fd_sc_hd__o22a_1
XFILLER_1_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_22_ _22_/A _22_/B VGND VGND VPWR VPWR _22_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_21_ _21_/A VGND VGND VPWR VPWR _21_/Y sky130_fd_sc_hd__inv_2
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_20_ _22_/A _22_/B _18_/Y _20_/B2 _19_/Y VGND VGND VPWR VPWR _21_/A sky130_fd_sc_hd__o221a_1
XFILLER_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput1 A_in[0] VGND VGND VPWR VPWR _24_/A sky130_fd_sc_hd__buf_1
XFILLER_10_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput2 A_in[1] VGND VGND VPWR VPWR _12_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 A_in[2] VGND VGND VPWR VPWR _20_/B2 sky130_fd_sc_hd__buf_1
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput4 A_in[3] VGND VGND VPWR VPWR _22_/A sky130_fd_sc_hd__buf_1
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput5 B_in[0] VGND VGND VPWR VPWR _13_/A sky130_fd_sc_hd__buf_1
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 B_in[1] VGND VGND VPWR VPWR _14_/A sky130_fd_sc_hd__buf_1
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
Xinput7 B_in[2] VGND VGND VPWR VPWR _18_/A sky130_fd_sc_hd__buf_1
XTAP_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput8 B_in[3] VGND VGND VPWR VPWR _17_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_22 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTAP_23 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_19_ _22_/A _22_/B _18_/Y _20_/B2 VGND VGND VPWR VPWR _19_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_24 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_18_ _18_/A VGND VGND VPWR VPWR _18_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_25 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_17_ _17_/A VGND VGND VPWR VPWR _22_/B sky130_fd_sc_hd__inv_2
XFILLER_5_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_26 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_16_ _14_/A _14_/B _15_/X VGND VGND VPWR VPWR _16_/X sky130_fd_sc_hd__o21ba_1
XFILLER_5_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_27 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_15_ _14_/A _14_/B _24_/A _13_/Y _14_/Y VGND VGND VPWR VPWR _15_/X sky130_fd_sc_hd__o221a_1
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_14_ _14_/A _14_/B VGND VGND VPWR VPWR _14_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_13_ _13_/A VGND VGND VPWR VPWR _13_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_5_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_12_ _12_/A VGND VGND VPWR VPWR _14_/B sky130_fd_sc_hd__inv_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_9_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
C163 _14_/B VGND 1.07fF
C164 _14_/Y VGND 1.46fF
C165 _13_/Y VGND 0.90fF
C166 _15_/X VGND 1.34fF
C167 _18_/Y VGND 0.35fF
C168 B_in[3] VGND 0.91fF
C169 _17_/A VGND 0.72fF
C170 B_in[2] VGND 0.77fF
C171 B_in[1] VGND 0.07fF
C172 B_in[0] VGND 0.84fF
C173 _13_/A VGND 1.55fF
C174 A_in[3] VGND 0.56fF
C175 A_in[2] VGND 0.79fF
C176 A_in[1] VGND 0.73fF
C177 A_in[0] VGND 0.85fF
C178 _19_/Y VGND 0.15fF
C179 _16_/X VGND 0.67fF
C180 _22_/Y VGND 1.05fF
C181 _21_/Y VGND 0.65fF
C182 _24_/Y VGND 1.35fF
C183 _26_/B VGND 3.22fF
C184 VPWR VGND 41.12fF
C185 less_than VGND 1.21fF
C186 equal_to VGND 0.81fF
C187 greater_than VGND 0.75fF
.ends
